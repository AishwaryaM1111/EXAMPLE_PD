magic
tech sky130A
magscale 1 2
timestamp 1740654827
<< nwell >>
rect 1066 2159 7398 8198
<< obsli1 >>
rect 1104 2159 7360 8177
<< obsm1 >>
rect 842 2128 7530 8208
<< obsm2 >>
rect 846 2139 7526 8197
<< metal3 >>
rect 0 5448 800 5568
rect 7735 5448 8535 5568
rect 0 4768 800 4888
rect 7735 4768 8535 4888
rect 0 4088 800 4208
<< obsm3 >>
rect 798 5648 7735 8193
rect 880 5368 7655 5648
rect 798 4968 7735 5368
rect 880 4688 7655 4968
rect 798 4288 7735 4688
rect 880 4008 7735 4288
rect 798 2143 7735 4008
<< metal4 >>
rect 1725 2128 2045 8208
rect 2385 2128 2705 8228
rect 3288 2128 3608 8208
rect 3948 2128 4268 8228
rect 4851 2128 5171 8208
rect 5511 2128 5831 8228
rect 6414 2128 6734 8208
rect 7074 2128 7394 8228
<< metal5 >>
rect 1056 7908 7408 8228
rect 1056 7248 7408 7568
rect 1056 6413 7408 6733
rect 1056 5753 7408 6073
rect 1056 4918 7408 5238
rect 1056 4258 7408 4578
rect 1056 3423 7408 3743
rect 1056 2763 7408 3083
<< labels >>
rlabel metal4 s 2385 2128 2705 8228 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3948 2128 4268 8228 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5511 2128 5831 8228 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7074 2128 7394 8228 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3423 7408 3743 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4918 7408 5238 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6413 7408 6733 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7908 7408 8228 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1725 2128 2045 8208 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3288 2128 3608 8208 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4851 2128 5171 8208 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6414 2128 6734 8208 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2763 7408 3083 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4258 7408 4578 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5753 7408 6073 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7248 7408 7568 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 5448 800 5568 6 a
port 3 nsew signal input
rlabel metal3 s 7735 4768 8535 4888 6 b
port 4 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 cin
port 5 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 co
port 6 nsew signal output
rlabel metal3 s 7735 5448 8535 5568 6 s
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 8535 10679
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 123064
string GDS_FILE /openlane/designs/new/runs/run1/results/signoff/new.magic.gds
string GDS_START 45866
<< end >>

