magic
tech sky130A
magscale 1 2
timestamp 1740654827
<< viali >>
rect 1409 5661 1443 5695
rect 6745 5661 6779 5695
rect 1593 5525 1627 5559
rect 6929 5525 6963 5559
rect 4445 5321 4479 5355
rect 3433 5253 3467 5287
rect 1685 5185 1719 5219
rect 3341 5185 3375 5219
rect 3617 5185 3651 5219
rect 4123 5185 4157 5219
rect 4905 5185 4939 5219
rect 7021 5185 7055 5219
rect 3985 5117 4019 5151
rect 4813 5117 4847 5151
rect 4537 5049 4571 5083
rect 6837 5049 6871 5083
rect 1501 4981 1535 5015
rect 3801 4981 3835 5015
rect 1593 4777 1627 4811
rect 3801 4777 3835 4811
rect 4169 4777 4203 4811
rect 4261 4641 4295 4675
rect 1409 4573 1443 4607
rect 3985 4573 4019 4607
<< metal1 >>
rect 1104 8186 7360 8208
rect 1104 8134 1731 8186
rect 1783 8134 1795 8186
rect 1847 8134 1859 8186
rect 1911 8134 1923 8186
rect 1975 8134 1987 8186
rect 2039 8134 3294 8186
rect 3346 8134 3358 8186
rect 3410 8134 3422 8186
rect 3474 8134 3486 8186
rect 3538 8134 3550 8186
rect 3602 8134 4857 8186
rect 4909 8134 4921 8186
rect 4973 8134 4985 8186
rect 5037 8134 5049 8186
rect 5101 8134 5113 8186
rect 5165 8134 6420 8186
rect 6472 8134 6484 8186
rect 6536 8134 6548 8186
rect 6600 8134 6612 8186
rect 6664 8134 6676 8186
rect 6728 8134 7360 8186
rect 1104 8112 7360 8134
rect 1104 7642 7394 7664
rect 1104 7590 2391 7642
rect 2443 7590 2455 7642
rect 2507 7590 2519 7642
rect 2571 7590 2583 7642
rect 2635 7590 2647 7642
rect 2699 7590 3954 7642
rect 4006 7590 4018 7642
rect 4070 7590 4082 7642
rect 4134 7590 4146 7642
rect 4198 7590 4210 7642
rect 4262 7590 5517 7642
rect 5569 7590 5581 7642
rect 5633 7590 5645 7642
rect 5697 7590 5709 7642
rect 5761 7590 5773 7642
rect 5825 7590 7080 7642
rect 7132 7590 7144 7642
rect 7196 7590 7208 7642
rect 7260 7590 7272 7642
rect 7324 7590 7336 7642
rect 7388 7590 7394 7642
rect 1104 7568 7394 7590
rect 1104 7098 7360 7120
rect 1104 7046 1731 7098
rect 1783 7046 1795 7098
rect 1847 7046 1859 7098
rect 1911 7046 1923 7098
rect 1975 7046 1987 7098
rect 2039 7046 3294 7098
rect 3346 7046 3358 7098
rect 3410 7046 3422 7098
rect 3474 7046 3486 7098
rect 3538 7046 3550 7098
rect 3602 7046 4857 7098
rect 4909 7046 4921 7098
rect 4973 7046 4985 7098
rect 5037 7046 5049 7098
rect 5101 7046 5113 7098
rect 5165 7046 6420 7098
rect 6472 7046 6484 7098
rect 6536 7046 6548 7098
rect 6600 7046 6612 7098
rect 6664 7046 6676 7098
rect 6728 7046 7360 7098
rect 1104 7024 7360 7046
rect 1104 6554 7394 6576
rect 1104 6502 2391 6554
rect 2443 6502 2455 6554
rect 2507 6502 2519 6554
rect 2571 6502 2583 6554
rect 2635 6502 2647 6554
rect 2699 6502 3954 6554
rect 4006 6502 4018 6554
rect 4070 6502 4082 6554
rect 4134 6502 4146 6554
rect 4198 6502 4210 6554
rect 4262 6502 5517 6554
rect 5569 6502 5581 6554
rect 5633 6502 5645 6554
rect 5697 6502 5709 6554
rect 5761 6502 5773 6554
rect 5825 6502 7080 6554
rect 7132 6502 7144 6554
rect 7196 6502 7208 6554
rect 7260 6502 7272 6554
rect 7324 6502 7336 6554
rect 7388 6502 7394 6554
rect 1104 6480 7394 6502
rect 1104 6010 7360 6032
rect 1104 5958 1731 6010
rect 1783 5958 1795 6010
rect 1847 5958 1859 6010
rect 1911 5958 1923 6010
rect 1975 5958 1987 6010
rect 2039 5958 3294 6010
rect 3346 5958 3358 6010
rect 3410 5958 3422 6010
rect 3474 5958 3486 6010
rect 3538 5958 3550 6010
rect 3602 5958 4857 6010
rect 4909 5958 4921 6010
rect 4973 5958 4985 6010
rect 5037 5958 5049 6010
rect 5101 5958 5113 6010
rect 5165 5958 6420 6010
rect 6472 5958 6484 6010
rect 6536 5958 6548 6010
rect 6600 5958 6612 6010
rect 6664 5958 6676 6010
rect 6728 5958 7360 6010
rect 1104 5936 7360 5958
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 6730 5652 6736 5704
rect 6788 5652 6794 5704
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 3326 5556 3332 5568
rect 1627 5528 3332 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 3326 5516 3332 5528
rect 3384 5556 3390 5568
rect 3878 5556 3884 5568
rect 3384 5528 3884 5556
rect 3384 5516 3390 5528
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7466 5556 7472 5568
rect 6963 5528 7472 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 1104 5466 7394 5488
rect 1104 5414 2391 5466
rect 2443 5414 2455 5466
rect 2507 5414 2519 5466
rect 2571 5414 2583 5466
rect 2635 5414 2647 5466
rect 2699 5414 3954 5466
rect 4006 5414 4018 5466
rect 4070 5414 4082 5466
rect 4134 5414 4146 5466
rect 4198 5414 4210 5466
rect 4262 5414 5517 5466
rect 5569 5414 5581 5466
rect 5633 5414 5645 5466
rect 5697 5414 5709 5466
rect 5761 5414 5773 5466
rect 5825 5414 7080 5466
rect 7132 5414 7144 5466
rect 7196 5414 7208 5466
rect 7260 5414 7272 5466
rect 7324 5414 7336 5466
rect 7388 5414 7394 5466
rect 1104 5392 7394 5414
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 6730 5352 6736 5364
rect 4479 5324 6736 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 3421 5287 3479 5293
rect 3421 5253 3433 5287
rect 3467 5284 3479 5287
rect 3467 5256 4936 5284
rect 3467 5253 3479 5256
rect 3421 5247 3479 5253
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 3142 5216 3148 5228
rect 1719 5188 3148 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 4908 5225 4936 5256
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 4111 5219 4169 5225
rect 4111 5216 4123 5219
rect 3651 5188 4123 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 4111 5185 4123 5188
rect 4157 5185 4169 5219
rect 4111 5179 4169 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 3620 5148 3648 5179
rect 1636 5120 3648 5148
rect 3973 5151 4031 5157
rect 1636 5108 1642 5120
rect 3973 5117 3985 5151
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 3988 5080 4016 5111
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4304 5120 4813 5148
rect 4304 5108 4310 5120
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 4525 5083 4583 5089
rect 4525 5080 4537 5083
rect 3988 5052 4537 5080
rect 4525 5049 4537 5052
rect 4571 5049 4583 5083
rect 4525 5043 4583 5049
rect 4614 5040 4620 5092
rect 4672 5080 4678 5092
rect 4908 5080 4936 5179
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 6825 5083 6883 5089
rect 6825 5080 6837 5083
rect 4672 5052 6837 5080
rect 4672 5040 4678 5052
rect 6825 5049 6837 5052
rect 6871 5049 6883 5083
rect 6825 5043 6883 5049
rect 842 4972 848 5024
rect 900 5012 906 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 900 4984 1501 5012
rect 900 4972 906 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 3789 5015 3847 5021
rect 3789 4981 3801 5015
rect 3835 5012 3847 5015
rect 3970 5012 3976 5024
rect 3835 4984 3976 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 1104 4922 7360 4944
rect 1104 4870 1731 4922
rect 1783 4870 1795 4922
rect 1847 4870 1859 4922
rect 1911 4870 1923 4922
rect 1975 4870 1987 4922
rect 2039 4870 3294 4922
rect 3346 4870 3358 4922
rect 3410 4870 3422 4922
rect 3474 4870 3486 4922
rect 3538 4870 3550 4922
rect 3602 4870 4857 4922
rect 4909 4870 4921 4922
rect 4973 4870 4985 4922
rect 5037 4870 5049 4922
rect 5101 4870 5113 4922
rect 5165 4870 6420 4922
rect 6472 4870 6484 4922
rect 6536 4870 6548 4922
rect 6600 4870 6612 4922
rect 6664 4870 6676 4922
rect 6728 4870 7360 4922
rect 1104 4848 7360 4870
rect 1578 4768 1584 4820
rect 1636 4768 1642 4820
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3200 4780 3801 4808
rect 3200 4768 3206 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 3936 4780 4169 4808
rect 3936 4768 3942 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4614 4672 4620 4684
rect 4295 4644 4620 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 1104 4378 7394 4400
rect 1104 4326 2391 4378
rect 2443 4326 2455 4378
rect 2507 4326 2519 4378
rect 2571 4326 2583 4378
rect 2635 4326 2647 4378
rect 2699 4326 3954 4378
rect 4006 4326 4018 4378
rect 4070 4326 4082 4378
rect 4134 4326 4146 4378
rect 4198 4326 4210 4378
rect 4262 4326 5517 4378
rect 5569 4326 5581 4378
rect 5633 4326 5645 4378
rect 5697 4326 5709 4378
rect 5761 4326 5773 4378
rect 5825 4326 7080 4378
rect 7132 4326 7144 4378
rect 7196 4326 7208 4378
rect 7260 4326 7272 4378
rect 7324 4326 7336 4378
rect 7388 4326 7394 4378
rect 1104 4304 7394 4326
rect 1104 3834 7360 3856
rect 1104 3782 1731 3834
rect 1783 3782 1795 3834
rect 1847 3782 1859 3834
rect 1911 3782 1923 3834
rect 1975 3782 1987 3834
rect 2039 3782 3294 3834
rect 3346 3782 3358 3834
rect 3410 3782 3422 3834
rect 3474 3782 3486 3834
rect 3538 3782 3550 3834
rect 3602 3782 4857 3834
rect 4909 3782 4921 3834
rect 4973 3782 4985 3834
rect 5037 3782 5049 3834
rect 5101 3782 5113 3834
rect 5165 3782 6420 3834
rect 6472 3782 6484 3834
rect 6536 3782 6548 3834
rect 6600 3782 6612 3834
rect 6664 3782 6676 3834
rect 6728 3782 7360 3834
rect 1104 3760 7360 3782
rect 1104 3290 7394 3312
rect 1104 3238 2391 3290
rect 2443 3238 2455 3290
rect 2507 3238 2519 3290
rect 2571 3238 2583 3290
rect 2635 3238 2647 3290
rect 2699 3238 3954 3290
rect 4006 3238 4018 3290
rect 4070 3238 4082 3290
rect 4134 3238 4146 3290
rect 4198 3238 4210 3290
rect 4262 3238 5517 3290
rect 5569 3238 5581 3290
rect 5633 3238 5645 3290
rect 5697 3238 5709 3290
rect 5761 3238 5773 3290
rect 5825 3238 7080 3290
rect 7132 3238 7144 3290
rect 7196 3238 7208 3290
rect 7260 3238 7272 3290
rect 7324 3238 7336 3290
rect 7388 3238 7394 3290
rect 1104 3216 7394 3238
rect 1104 2746 7360 2768
rect 1104 2694 1731 2746
rect 1783 2694 1795 2746
rect 1847 2694 1859 2746
rect 1911 2694 1923 2746
rect 1975 2694 1987 2746
rect 2039 2694 3294 2746
rect 3346 2694 3358 2746
rect 3410 2694 3422 2746
rect 3474 2694 3486 2746
rect 3538 2694 3550 2746
rect 3602 2694 4857 2746
rect 4909 2694 4921 2746
rect 4973 2694 4985 2746
rect 5037 2694 5049 2746
rect 5101 2694 5113 2746
rect 5165 2694 6420 2746
rect 6472 2694 6484 2746
rect 6536 2694 6548 2746
rect 6600 2694 6612 2746
rect 6664 2694 6676 2746
rect 6728 2694 7360 2746
rect 1104 2672 7360 2694
rect 1104 2202 7394 2224
rect 1104 2150 2391 2202
rect 2443 2150 2455 2202
rect 2507 2150 2519 2202
rect 2571 2150 2583 2202
rect 2635 2150 2647 2202
rect 2699 2150 3954 2202
rect 4006 2150 4018 2202
rect 4070 2150 4082 2202
rect 4134 2150 4146 2202
rect 4198 2150 4210 2202
rect 4262 2150 5517 2202
rect 5569 2150 5581 2202
rect 5633 2150 5645 2202
rect 5697 2150 5709 2202
rect 5761 2150 5773 2202
rect 5825 2150 7080 2202
rect 7132 2150 7144 2202
rect 7196 2150 7208 2202
rect 7260 2150 7272 2202
rect 7324 2150 7336 2202
rect 7388 2150 7394 2202
rect 1104 2128 7394 2150
<< via1 >>
rect 1731 8134 1783 8186
rect 1795 8134 1847 8186
rect 1859 8134 1911 8186
rect 1923 8134 1975 8186
rect 1987 8134 2039 8186
rect 3294 8134 3346 8186
rect 3358 8134 3410 8186
rect 3422 8134 3474 8186
rect 3486 8134 3538 8186
rect 3550 8134 3602 8186
rect 4857 8134 4909 8186
rect 4921 8134 4973 8186
rect 4985 8134 5037 8186
rect 5049 8134 5101 8186
rect 5113 8134 5165 8186
rect 6420 8134 6472 8186
rect 6484 8134 6536 8186
rect 6548 8134 6600 8186
rect 6612 8134 6664 8186
rect 6676 8134 6728 8186
rect 2391 7590 2443 7642
rect 2455 7590 2507 7642
rect 2519 7590 2571 7642
rect 2583 7590 2635 7642
rect 2647 7590 2699 7642
rect 3954 7590 4006 7642
rect 4018 7590 4070 7642
rect 4082 7590 4134 7642
rect 4146 7590 4198 7642
rect 4210 7590 4262 7642
rect 5517 7590 5569 7642
rect 5581 7590 5633 7642
rect 5645 7590 5697 7642
rect 5709 7590 5761 7642
rect 5773 7590 5825 7642
rect 7080 7590 7132 7642
rect 7144 7590 7196 7642
rect 7208 7590 7260 7642
rect 7272 7590 7324 7642
rect 7336 7590 7388 7642
rect 1731 7046 1783 7098
rect 1795 7046 1847 7098
rect 1859 7046 1911 7098
rect 1923 7046 1975 7098
rect 1987 7046 2039 7098
rect 3294 7046 3346 7098
rect 3358 7046 3410 7098
rect 3422 7046 3474 7098
rect 3486 7046 3538 7098
rect 3550 7046 3602 7098
rect 4857 7046 4909 7098
rect 4921 7046 4973 7098
rect 4985 7046 5037 7098
rect 5049 7046 5101 7098
rect 5113 7046 5165 7098
rect 6420 7046 6472 7098
rect 6484 7046 6536 7098
rect 6548 7046 6600 7098
rect 6612 7046 6664 7098
rect 6676 7046 6728 7098
rect 2391 6502 2443 6554
rect 2455 6502 2507 6554
rect 2519 6502 2571 6554
rect 2583 6502 2635 6554
rect 2647 6502 2699 6554
rect 3954 6502 4006 6554
rect 4018 6502 4070 6554
rect 4082 6502 4134 6554
rect 4146 6502 4198 6554
rect 4210 6502 4262 6554
rect 5517 6502 5569 6554
rect 5581 6502 5633 6554
rect 5645 6502 5697 6554
rect 5709 6502 5761 6554
rect 5773 6502 5825 6554
rect 7080 6502 7132 6554
rect 7144 6502 7196 6554
rect 7208 6502 7260 6554
rect 7272 6502 7324 6554
rect 7336 6502 7388 6554
rect 1731 5958 1783 6010
rect 1795 5958 1847 6010
rect 1859 5958 1911 6010
rect 1923 5958 1975 6010
rect 1987 5958 2039 6010
rect 3294 5958 3346 6010
rect 3358 5958 3410 6010
rect 3422 5958 3474 6010
rect 3486 5958 3538 6010
rect 3550 5958 3602 6010
rect 4857 5958 4909 6010
rect 4921 5958 4973 6010
rect 4985 5958 5037 6010
rect 5049 5958 5101 6010
rect 5113 5958 5165 6010
rect 6420 5958 6472 6010
rect 6484 5958 6536 6010
rect 6548 5958 6600 6010
rect 6612 5958 6664 6010
rect 6676 5958 6728 6010
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 6736 5695 6788 5704
rect 6736 5661 6745 5695
rect 6745 5661 6779 5695
rect 6779 5661 6788 5695
rect 6736 5652 6788 5661
rect 3332 5516 3384 5568
rect 3884 5516 3936 5568
rect 7472 5516 7524 5568
rect 2391 5414 2443 5466
rect 2455 5414 2507 5466
rect 2519 5414 2571 5466
rect 2583 5414 2635 5466
rect 2647 5414 2699 5466
rect 3954 5414 4006 5466
rect 4018 5414 4070 5466
rect 4082 5414 4134 5466
rect 4146 5414 4198 5466
rect 4210 5414 4262 5466
rect 5517 5414 5569 5466
rect 5581 5414 5633 5466
rect 5645 5414 5697 5466
rect 5709 5414 5761 5466
rect 5773 5414 5825 5466
rect 7080 5414 7132 5466
rect 7144 5414 7196 5466
rect 7208 5414 7260 5466
rect 7272 5414 7324 5466
rect 7336 5414 7388 5466
rect 6736 5312 6788 5364
rect 3148 5176 3200 5228
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 1584 5108 1636 5160
rect 4252 5108 4304 5160
rect 4620 5040 4672 5092
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 848 4972 900 5024
rect 3976 4972 4028 5024
rect 1731 4870 1783 4922
rect 1795 4870 1847 4922
rect 1859 4870 1911 4922
rect 1923 4870 1975 4922
rect 1987 4870 2039 4922
rect 3294 4870 3346 4922
rect 3358 4870 3410 4922
rect 3422 4870 3474 4922
rect 3486 4870 3538 4922
rect 3550 4870 3602 4922
rect 4857 4870 4909 4922
rect 4921 4870 4973 4922
rect 4985 4870 5037 4922
rect 5049 4870 5101 4922
rect 5113 4870 5165 4922
rect 6420 4870 6472 4922
rect 6484 4870 6536 4922
rect 6548 4870 6600 4922
rect 6612 4870 6664 4922
rect 6676 4870 6728 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 3148 4768 3200 4820
rect 3884 4768 3936 4820
rect 4620 4632 4672 4684
rect 848 4564 900 4616
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 2391 4326 2443 4378
rect 2455 4326 2507 4378
rect 2519 4326 2571 4378
rect 2583 4326 2635 4378
rect 2647 4326 2699 4378
rect 3954 4326 4006 4378
rect 4018 4326 4070 4378
rect 4082 4326 4134 4378
rect 4146 4326 4198 4378
rect 4210 4326 4262 4378
rect 5517 4326 5569 4378
rect 5581 4326 5633 4378
rect 5645 4326 5697 4378
rect 5709 4326 5761 4378
rect 5773 4326 5825 4378
rect 7080 4326 7132 4378
rect 7144 4326 7196 4378
rect 7208 4326 7260 4378
rect 7272 4326 7324 4378
rect 7336 4326 7388 4378
rect 1731 3782 1783 3834
rect 1795 3782 1847 3834
rect 1859 3782 1911 3834
rect 1923 3782 1975 3834
rect 1987 3782 2039 3834
rect 3294 3782 3346 3834
rect 3358 3782 3410 3834
rect 3422 3782 3474 3834
rect 3486 3782 3538 3834
rect 3550 3782 3602 3834
rect 4857 3782 4909 3834
rect 4921 3782 4973 3834
rect 4985 3782 5037 3834
rect 5049 3782 5101 3834
rect 5113 3782 5165 3834
rect 6420 3782 6472 3834
rect 6484 3782 6536 3834
rect 6548 3782 6600 3834
rect 6612 3782 6664 3834
rect 6676 3782 6728 3834
rect 2391 3238 2443 3290
rect 2455 3238 2507 3290
rect 2519 3238 2571 3290
rect 2583 3238 2635 3290
rect 2647 3238 2699 3290
rect 3954 3238 4006 3290
rect 4018 3238 4070 3290
rect 4082 3238 4134 3290
rect 4146 3238 4198 3290
rect 4210 3238 4262 3290
rect 5517 3238 5569 3290
rect 5581 3238 5633 3290
rect 5645 3238 5697 3290
rect 5709 3238 5761 3290
rect 5773 3238 5825 3290
rect 7080 3238 7132 3290
rect 7144 3238 7196 3290
rect 7208 3238 7260 3290
rect 7272 3238 7324 3290
rect 7336 3238 7388 3290
rect 1731 2694 1783 2746
rect 1795 2694 1847 2746
rect 1859 2694 1911 2746
rect 1923 2694 1975 2746
rect 1987 2694 2039 2746
rect 3294 2694 3346 2746
rect 3358 2694 3410 2746
rect 3422 2694 3474 2746
rect 3486 2694 3538 2746
rect 3550 2694 3602 2746
rect 4857 2694 4909 2746
rect 4921 2694 4973 2746
rect 4985 2694 5037 2746
rect 5049 2694 5101 2746
rect 5113 2694 5165 2746
rect 6420 2694 6472 2746
rect 6484 2694 6536 2746
rect 6548 2694 6600 2746
rect 6612 2694 6664 2746
rect 6676 2694 6728 2746
rect 2391 2150 2443 2202
rect 2455 2150 2507 2202
rect 2519 2150 2571 2202
rect 2583 2150 2635 2202
rect 2647 2150 2699 2202
rect 3954 2150 4006 2202
rect 4018 2150 4070 2202
rect 4082 2150 4134 2202
rect 4146 2150 4198 2202
rect 4210 2150 4262 2202
rect 5517 2150 5569 2202
rect 5581 2150 5633 2202
rect 5645 2150 5697 2202
rect 5709 2150 5761 2202
rect 5773 2150 5825 2202
rect 7080 2150 7132 2202
rect 7144 2150 7196 2202
rect 7208 2150 7260 2202
rect 7272 2150 7324 2202
rect 7336 2150 7388 2202
<< metal2 >>
rect 1731 8188 2039 8197
rect 1731 8186 1737 8188
rect 1793 8186 1817 8188
rect 1873 8186 1897 8188
rect 1953 8186 1977 8188
rect 2033 8186 2039 8188
rect 1793 8134 1795 8186
rect 1975 8134 1977 8186
rect 1731 8132 1737 8134
rect 1793 8132 1817 8134
rect 1873 8132 1897 8134
rect 1953 8132 1977 8134
rect 2033 8132 2039 8134
rect 1731 8123 2039 8132
rect 3294 8188 3602 8197
rect 3294 8186 3300 8188
rect 3356 8186 3380 8188
rect 3436 8186 3460 8188
rect 3516 8186 3540 8188
rect 3596 8186 3602 8188
rect 3356 8134 3358 8186
rect 3538 8134 3540 8186
rect 3294 8132 3300 8134
rect 3356 8132 3380 8134
rect 3436 8132 3460 8134
rect 3516 8132 3540 8134
rect 3596 8132 3602 8134
rect 3294 8123 3602 8132
rect 4857 8188 5165 8197
rect 4857 8186 4863 8188
rect 4919 8186 4943 8188
rect 4999 8186 5023 8188
rect 5079 8186 5103 8188
rect 5159 8186 5165 8188
rect 4919 8134 4921 8186
rect 5101 8134 5103 8186
rect 4857 8132 4863 8134
rect 4919 8132 4943 8134
rect 4999 8132 5023 8134
rect 5079 8132 5103 8134
rect 5159 8132 5165 8134
rect 4857 8123 5165 8132
rect 6420 8188 6728 8197
rect 6420 8186 6426 8188
rect 6482 8186 6506 8188
rect 6562 8186 6586 8188
rect 6642 8186 6666 8188
rect 6722 8186 6728 8188
rect 6482 8134 6484 8186
rect 6664 8134 6666 8186
rect 6420 8132 6426 8134
rect 6482 8132 6506 8134
rect 6562 8132 6586 8134
rect 6642 8132 6666 8134
rect 6722 8132 6728 8134
rect 6420 8123 6728 8132
rect 2391 7644 2699 7653
rect 2391 7642 2397 7644
rect 2453 7642 2477 7644
rect 2533 7642 2557 7644
rect 2613 7642 2637 7644
rect 2693 7642 2699 7644
rect 2453 7590 2455 7642
rect 2635 7590 2637 7642
rect 2391 7588 2397 7590
rect 2453 7588 2477 7590
rect 2533 7588 2557 7590
rect 2613 7588 2637 7590
rect 2693 7588 2699 7590
rect 2391 7579 2699 7588
rect 3954 7644 4262 7653
rect 3954 7642 3960 7644
rect 4016 7642 4040 7644
rect 4096 7642 4120 7644
rect 4176 7642 4200 7644
rect 4256 7642 4262 7644
rect 4016 7590 4018 7642
rect 4198 7590 4200 7642
rect 3954 7588 3960 7590
rect 4016 7588 4040 7590
rect 4096 7588 4120 7590
rect 4176 7588 4200 7590
rect 4256 7588 4262 7590
rect 3954 7579 4262 7588
rect 5517 7644 5825 7653
rect 5517 7642 5523 7644
rect 5579 7642 5603 7644
rect 5659 7642 5683 7644
rect 5739 7642 5763 7644
rect 5819 7642 5825 7644
rect 5579 7590 5581 7642
rect 5761 7590 5763 7642
rect 5517 7588 5523 7590
rect 5579 7588 5603 7590
rect 5659 7588 5683 7590
rect 5739 7588 5763 7590
rect 5819 7588 5825 7590
rect 5517 7579 5825 7588
rect 7080 7644 7388 7653
rect 7080 7642 7086 7644
rect 7142 7642 7166 7644
rect 7222 7642 7246 7644
rect 7302 7642 7326 7644
rect 7382 7642 7388 7644
rect 7142 7590 7144 7642
rect 7324 7590 7326 7642
rect 7080 7588 7086 7590
rect 7142 7588 7166 7590
rect 7222 7588 7246 7590
rect 7302 7588 7326 7590
rect 7382 7588 7388 7590
rect 7080 7579 7388 7588
rect 1731 7100 2039 7109
rect 1731 7098 1737 7100
rect 1793 7098 1817 7100
rect 1873 7098 1897 7100
rect 1953 7098 1977 7100
rect 2033 7098 2039 7100
rect 1793 7046 1795 7098
rect 1975 7046 1977 7098
rect 1731 7044 1737 7046
rect 1793 7044 1817 7046
rect 1873 7044 1897 7046
rect 1953 7044 1977 7046
rect 2033 7044 2039 7046
rect 1731 7035 2039 7044
rect 3294 7100 3602 7109
rect 3294 7098 3300 7100
rect 3356 7098 3380 7100
rect 3436 7098 3460 7100
rect 3516 7098 3540 7100
rect 3596 7098 3602 7100
rect 3356 7046 3358 7098
rect 3538 7046 3540 7098
rect 3294 7044 3300 7046
rect 3356 7044 3380 7046
rect 3436 7044 3460 7046
rect 3516 7044 3540 7046
rect 3596 7044 3602 7046
rect 3294 7035 3602 7044
rect 4857 7100 5165 7109
rect 4857 7098 4863 7100
rect 4919 7098 4943 7100
rect 4999 7098 5023 7100
rect 5079 7098 5103 7100
rect 5159 7098 5165 7100
rect 4919 7046 4921 7098
rect 5101 7046 5103 7098
rect 4857 7044 4863 7046
rect 4919 7044 4943 7046
rect 4999 7044 5023 7046
rect 5079 7044 5103 7046
rect 5159 7044 5165 7046
rect 4857 7035 5165 7044
rect 6420 7100 6728 7109
rect 6420 7098 6426 7100
rect 6482 7098 6506 7100
rect 6562 7098 6586 7100
rect 6642 7098 6666 7100
rect 6722 7098 6728 7100
rect 6482 7046 6484 7098
rect 6664 7046 6666 7098
rect 6420 7044 6426 7046
rect 6482 7044 6506 7046
rect 6562 7044 6586 7046
rect 6642 7044 6666 7046
rect 6722 7044 6728 7046
rect 6420 7035 6728 7044
rect 2391 6556 2699 6565
rect 2391 6554 2397 6556
rect 2453 6554 2477 6556
rect 2533 6554 2557 6556
rect 2613 6554 2637 6556
rect 2693 6554 2699 6556
rect 2453 6502 2455 6554
rect 2635 6502 2637 6554
rect 2391 6500 2397 6502
rect 2453 6500 2477 6502
rect 2533 6500 2557 6502
rect 2613 6500 2637 6502
rect 2693 6500 2699 6502
rect 2391 6491 2699 6500
rect 3954 6556 4262 6565
rect 3954 6554 3960 6556
rect 4016 6554 4040 6556
rect 4096 6554 4120 6556
rect 4176 6554 4200 6556
rect 4256 6554 4262 6556
rect 4016 6502 4018 6554
rect 4198 6502 4200 6554
rect 3954 6500 3960 6502
rect 4016 6500 4040 6502
rect 4096 6500 4120 6502
rect 4176 6500 4200 6502
rect 4256 6500 4262 6502
rect 3954 6491 4262 6500
rect 5517 6556 5825 6565
rect 5517 6554 5523 6556
rect 5579 6554 5603 6556
rect 5659 6554 5683 6556
rect 5739 6554 5763 6556
rect 5819 6554 5825 6556
rect 5579 6502 5581 6554
rect 5761 6502 5763 6554
rect 5517 6500 5523 6502
rect 5579 6500 5603 6502
rect 5659 6500 5683 6502
rect 5739 6500 5763 6502
rect 5819 6500 5825 6502
rect 5517 6491 5825 6500
rect 7080 6556 7388 6565
rect 7080 6554 7086 6556
rect 7142 6554 7166 6556
rect 7222 6554 7246 6556
rect 7302 6554 7326 6556
rect 7382 6554 7388 6556
rect 7142 6502 7144 6554
rect 7324 6502 7326 6554
rect 7080 6500 7086 6502
rect 7142 6500 7166 6502
rect 7222 6500 7246 6502
rect 7302 6500 7326 6502
rect 7382 6500 7388 6502
rect 7080 6491 7388 6500
rect 1731 6012 2039 6021
rect 1731 6010 1737 6012
rect 1793 6010 1817 6012
rect 1873 6010 1897 6012
rect 1953 6010 1977 6012
rect 2033 6010 2039 6012
rect 1793 5958 1795 6010
rect 1975 5958 1977 6010
rect 1731 5956 1737 5958
rect 1793 5956 1817 5958
rect 1873 5956 1897 5958
rect 1953 5956 1977 5958
rect 2033 5956 2039 5958
rect 1731 5947 2039 5956
rect 3294 6012 3602 6021
rect 3294 6010 3300 6012
rect 3356 6010 3380 6012
rect 3436 6010 3460 6012
rect 3516 6010 3540 6012
rect 3596 6010 3602 6012
rect 3356 5958 3358 6010
rect 3538 5958 3540 6010
rect 3294 5956 3300 5958
rect 3356 5956 3380 5958
rect 3436 5956 3460 5958
rect 3516 5956 3540 5958
rect 3596 5956 3602 5958
rect 3294 5947 3602 5956
rect 4857 6012 5165 6021
rect 4857 6010 4863 6012
rect 4919 6010 4943 6012
rect 4999 6010 5023 6012
rect 5079 6010 5103 6012
rect 5159 6010 5165 6012
rect 4919 5958 4921 6010
rect 5101 5958 5103 6010
rect 4857 5956 4863 5958
rect 4919 5956 4943 5958
rect 4999 5956 5023 5958
rect 5079 5956 5103 5958
rect 5159 5956 5165 5958
rect 4857 5947 5165 5956
rect 6420 6012 6728 6021
rect 6420 6010 6426 6012
rect 6482 6010 6506 6012
rect 6562 6010 6586 6012
rect 6642 6010 6666 6012
rect 6722 6010 6728 6012
rect 6482 5958 6484 6010
rect 6664 5958 6666 6010
rect 6420 5956 6426 5958
rect 6482 5956 6506 5958
rect 6562 5956 6586 5958
rect 6642 5956 6666 5958
rect 6722 5956 6728 5958
rect 6420 5947 6728 5956
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 1412 5545 1440 5646
rect 3332 5568 3384 5574
rect 1398 5536 1454 5545
rect 3332 5510 3384 5516
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 1398 5471 1454 5480
rect 2391 5468 2699 5477
rect 2391 5466 2397 5468
rect 2453 5466 2477 5468
rect 2533 5466 2557 5468
rect 2613 5466 2637 5468
rect 2693 5466 2699 5468
rect 2453 5414 2455 5466
rect 2635 5414 2637 5466
rect 2391 5412 2397 5414
rect 2453 5412 2477 5414
rect 2533 5412 2557 5414
rect 2613 5412 2637 5414
rect 2693 5412 2699 5414
rect 2391 5403 2699 5412
rect 3344 5234 3372 5510
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 848 5024 900 5030
rect 846 4992 848 5001
rect 900 4992 902 5001
rect 846 4927 902 4936
rect 1596 4826 1624 5102
rect 1731 4924 2039 4933
rect 1731 4922 1737 4924
rect 1793 4922 1817 4924
rect 1873 4922 1897 4924
rect 1953 4922 1977 4924
rect 2033 4922 2039 4924
rect 1793 4870 1795 4922
rect 1975 4870 1977 4922
rect 1731 4868 1737 4870
rect 1793 4868 1817 4870
rect 1873 4868 1897 4870
rect 1953 4868 1977 4870
rect 2033 4868 2039 4870
rect 1731 4859 2039 4868
rect 3160 4826 3188 5170
rect 3896 5114 3924 5510
rect 3954 5468 4262 5477
rect 3954 5466 3960 5468
rect 4016 5466 4040 5468
rect 4096 5466 4120 5468
rect 4176 5466 4200 5468
rect 4256 5466 4262 5468
rect 4016 5414 4018 5466
rect 4198 5414 4200 5466
rect 3954 5412 3960 5414
rect 4016 5412 4040 5414
rect 4096 5412 4120 5414
rect 4176 5412 4200 5414
rect 4256 5412 4262 5414
rect 3954 5403 4262 5412
rect 5517 5468 5825 5477
rect 5517 5466 5523 5468
rect 5579 5466 5603 5468
rect 5659 5466 5683 5468
rect 5739 5466 5763 5468
rect 5819 5466 5825 5468
rect 5579 5414 5581 5466
rect 5761 5414 5763 5466
rect 5517 5412 5523 5414
rect 5579 5412 5603 5414
rect 5659 5412 5683 5414
rect 5739 5412 5763 5414
rect 5819 5412 5825 5414
rect 5517 5403 5825 5412
rect 6748 5370 6776 5646
rect 7472 5568 7524 5574
rect 7470 5536 7472 5545
rect 7524 5536 7526 5545
rect 7080 5468 7388 5477
rect 7470 5471 7526 5480
rect 7080 5466 7086 5468
rect 7142 5466 7166 5468
rect 7222 5466 7246 5468
rect 7302 5466 7326 5468
rect 7382 5466 7388 5468
rect 7142 5414 7144 5466
rect 7324 5414 7326 5466
rect 7080 5412 7086 5414
rect 7142 5412 7166 5414
rect 7222 5412 7246 5414
rect 7302 5412 7326 5414
rect 7382 5412 7388 5414
rect 7080 5403 7388 5412
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 4252 5160 4304 5166
rect 3896 5108 4252 5114
rect 3896 5102 4304 5108
rect 3896 5086 4292 5102
rect 4620 5092 4672 5098
rect 3294 4924 3602 4933
rect 3294 4922 3300 4924
rect 3356 4922 3380 4924
rect 3436 4922 3460 4924
rect 3516 4922 3540 4924
rect 3596 4922 3602 4924
rect 3356 4870 3358 4922
rect 3538 4870 3540 4922
rect 3294 4868 3300 4870
rect 3356 4868 3380 4870
rect 3436 4868 3460 4870
rect 3516 4868 3540 4870
rect 3596 4868 3602 4870
rect 3294 4859 3602 4868
rect 3896 4826 3924 5086
rect 4620 5034 4672 5040
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3988 4622 4016 4966
rect 4632 4690 4660 5034
rect 4857 4924 5165 4933
rect 4857 4922 4863 4924
rect 4919 4922 4943 4924
rect 4999 4922 5023 4924
rect 5079 4922 5103 4924
rect 5159 4922 5165 4924
rect 4919 4870 4921 4922
rect 5101 4870 5103 4922
rect 4857 4868 4863 4870
rect 4919 4868 4943 4870
rect 4999 4868 5023 4870
rect 5079 4868 5103 4870
rect 5159 4868 5165 4870
rect 4857 4859 5165 4868
rect 6420 4924 6728 4933
rect 6420 4922 6426 4924
rect 6482 4922 6506 4924
rect 6562 4922 6586 4924
rect 6642 4922 6666 4924
rect 6722 4922 6728 4924
rect 6482 4870 6484 4922
rect 6664 4870 6666 4922
rect 6420 4868 6426 4870
rect 6482 4868 6506 4870
rect 6562 4868 6586 4870
rect 6642 4868 6666 4870
rect 6722 4868 6728 4870
rect 6420 4859 6728 4868
rect 7024 4865 7052 5170
rect 7010 4856 7066 4865
rect 7010 4791 7066 4800
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 860 4321 888 4558
rect 2391 4380 2699 4389
rect 2391 4378 2397 4380
rect 2453 4378 2477 4380
rect 2533 4378 2557 4380
rect 2613 4378 2637 4380
rect 2693 4378 2699 4380
rect 2453 4326 2455 4378
rect 2635 4326 2637 4378
rect 2391 4324 2397 4326
rect 2453 4324 2477 4326
rect 2533 4324 2557 4326
rect 2613 4324 2637 4326
rect 2693 4324 2699 4326
rect 846 4312 902 4321
rect 2391 4315 2699 4324
rect 3954 4380 4262 4389
rect 3954 4378 3960 4380
rect 4016 4378 4040 4380
rect 4096 4378 4120 4380
rect 4176 4378 4200 4380
rect 4256 4378 4262 4380
rect 4016 4326 4018 4378
rect 4198 4326 4200 4378
rect 3954 4324 3960 4326
rect 4016 4324 4040 4326
rect 4096 4324 4120 4326
rect 4176 4324 4200 4326
rect 4256 4324 4262 4326
rect 3954 4315 4262 4324
rect 5517 4380 5825 4389
rect 5517 4378 5523 4380
rect 5579 4378 5603 4380
rect 5659 4378 5683 4380
rect 5739 4378 5763 4380
rect 5819 4378 5825 4380
rect 5579 4326 5581 4378
rect 5761 4326 5763 4378
rect 5517 4324 5523 4326
rect 5579 4324 5603 4326
rect 5659 4324 5683 4326
rect 5739 4324 5763 4326
rect 5819 4324 5825 4326
rect 5517 4315 5825 4324
rect 7080 4380 7388 4389
rect 7080 4378 7086 4380
rect 7142 4378 7166 4380
rect 7222 4378 7246 4380
rect 7302 4378 7326 4380
rect 7382 4378 7388 4380
rect 7142 4326 7144 4378
rect 7324 4326 7326 4378
rect 7080 4324 7086 4326
rect 7142 4324 7166 4326
rect 7222 4324 7246 4326
rect 7302 4324 7326 4326
rect 7382 4324 7388 4326
rect 7080 4315 7388 4324
rect 846 4247 902 4256
rect 1731 3836 2039 3845
rect 1731 3834 1737 3836
rect 1793 3834 1817 3836
rect 1873 3834 1897 3836
rect 1953 3834 1977 3836
rect 2033 3834 2039 3836
rect 1793 3782 1795 3834
rect 1975 3782 1977 3834
rect 1731 3780 1737 3782
rect 1793 3780 1817 3782
rect 1873 3780 1897 3782
rect 1953 3780 1977 3782
rect 2033 3780 2039 3782
rect 1731 3771 2039 3780
rect 3294 3836 3602 3845
rect 3294 3834 3300 3836
rect 3356 3834 3380 3836
rect 3436 3834 3460 3836
rect 3516 3834 3540 3836
rect 3596 3834 3602 3836
rect 3356 3782 3358 3834
rect 3538 3782 3540 3834
rect 3294 3780 3300 3782
rect 3356 3780 3380 3782
rect 3436 3780 3460 3782
rect 3516 3780 3540 3782
rect 3596 3780 3602 3782
rect 3294 3771 3602 3780
rect 4857 3836 5165 3845
rect 4857 3834 4863 3836
rect 4919 3834 4943 3836
rect 4999 3834 5023 3836
rect 5079 3834 5103 3836
rect 5159 3834 5165 3836
rect 4919 3782 4921 3834
rect 5101 3782 5103 3834
rect 4857 3780 4863 3782
rect 4919 3780 4943 3782
rect 4999 3780 5023 3782
rect 5079 3780 5103 3782
rect 5159 3780 5165 3782
rect 4857 3771 5165 3780
rect 6420 3836 6728 3845
rect 6420 3834 6426 3836
rect 6482 3834 6506 3836
rect 6562 3834 6586 3836
rect 6642 3834 6666 3836
rect 6722 3834 6728 3836
rect 6482 3782 6484 3834
rect 6664 3782 6666 3834
rect 6420 3780 6426 3782
rect 6482 3780 6506 3782
rect 6562 3780 6586 3782
rect 6642 3780 6666 3782
rect 6722 3780 6728 3782
rect 6420 3771 6728 3780
rect 2391 3292 2699 3301
rect 2391 3290 2397 3292
rect 2453 3290 2477 3292
rect 2533 3290 2557 3292
rect 2613 3290 2637 3292
rect 2693 3290 2699 3292
rect 2453 3238 2455 3290
rect 2635 3238 2637 3290
rect 2391 3236 2397 3238
rect 2453 3236 2477 3238
rect 2533 3236 2557 3238
rect 2613 3236 2637 3238
rect 2693 3236 2699 3238
rect 2391 3227 2699 3236
rect 3954 3292 4262 3301
rect 3954 3290 3960 3292
rect 4016 3290 4040 3292
rect 4096 3290 4120 3292
rect 4176 3290 4200 3292
rect 4256 3290 4262 3292
rect 4016 3238 4018 3290
rect 4198 3238 4200 3290
rect 3954 3236 3960 3238
rect 4016 3236 4040 3238
rect 4096 3236 4120 3238
rect 4176 3236 4200 3238
rect 4256 3236 4262 3238
rect 3954 3227 4262 3236
rect 5517 3292 5825 3301
rect 5517 3290 5523 3292
rect 5579 3290 5603 3292
rect 5659 3290 5683 3292
rect 5739 3290 5763 3292
rect 5819 3290 5825 3292
rect 5579 3238 5581 3290
rect 5761 3238 5763 3290
rect 5517 3236 5523 3238
rect 5579 3236 5603 3238
rect 5659 3236 5683 3238
rect 5739 3236 5763 3238
rect 5819 3236 5825 3238
rect 5517 3227 5825 3236
rect 7080 3292 7388 3301
rect 7080 3290 7086 3292
rect 7142 3290 7166 3292
rect 7222 3290 7246 3292
rect 7302 3290 7326 3292
rect 7382 3290 7388 3292
rect 7142 3238 7144 3290
rect 7324 3238 7326 3290
rect 7080 3236 7086 3238
rect 7142 3236 7166 3238
rect 7222 3236 7246 3238
rect 7302 3236 7326 3238
rect 7382 3236 7388 3238
rect 7080 3227 7388 3236
rect 1731 2748 2039 2757
rect 1731 2746 1737 2748
rect 1793 2746 1817 2748
rect 1873 2746 1897 2748
rect 1953 2746 1977 2748
rect 2033 2746 2039 2748
rect 1793 2694 1795 2746
rect 1975 2694 1977 2746
rect 1731 2692 1737 2694
rect 1793 2692 1817 2694
rect 1873 2692 1897 2694
rect 1953 2692 1977 2694
rect 2033 2692 2039 2694
rect 1731 2683 2039 2692
rect 3294 2748 3602 2757
rect 3294 2746 3300 2748
rect 3356 2746 3380 2748
rect 3436 2746 3460 2748
rect 3516 2746 3540 2748
rect 3596 2746 3602 2748
rect 3356 2694 3358 2746
rect 3538 2694 3540 2746
rect 3294 2692 3300 2694
rect 3356 2692 3380 2694
rect 3436 2692 3460 2694
rect 3516 2692 3540 2694
rect 3596 2692 3602 2694
rect 3294 2683 3602 2692
rect 4857 2748 5165 2757
rect 4857 2746 4863 2748
rect 4919 2746 4943 2748
rect 4999 2746 5023 2748
rect 5079 2746 5103 2748
rect 5159 2746 5165 2748
rect 4919 2694 4921 2746
rect 5101 2694 5103 2746
rect 4857 2692 4863 2694
rect 4919 2692 4943 2694
rect 4999 2692 5023 2694
rect 5079 2692 5103 2694
rect 5159 2692 5165 2694
rect 4857 2683 5165 2692
rect 6420 2748 6728 2757
rect 6420 2746 6426 2748
rect 6482 2746 6506 2748
rect 6562 2746 6586 2748
rect 6642 2746 6666 2748
rect 6722 2746 6728 2748
rect 6482 2694 6484 2746
rect 6664 2694 6666 2746
rect 6420 2692 6426 2694
rect 6482 2692 6506 2694
rect 6562 2692 6586 2694
rect 6642 2692 6666 2694
rect 6722 2692 6728 2694
rect 6420 2683 6728 2692
rect 2391 2204 2699 2213
rect 2391 2202 2397 2204
rect 2453 2202 2477 2204
rect 2533 2202 2557 2204
rect 2613 2202 2637 2204
rect 2693 2202 2699 2204
rect 2453 2150 2455 2202
rect 2635 2150 2637 2202
rect 2391 2148 2397 2150
rect 2453 2148 2477 2150
rect 2533 2148 2557 2150
rect 2613 2148 2637 2150
rect 2693 2148 2699 2150
rect 2391 2139 2699 2148
rect 3954 2204 4262 2213
rect 3954 2202 3960 2204
rect 4016 2202 4040 2204
rect 4096 2202 4120 2204
rect 4176 2202 4200 2204
rect 4256 2202 4262 2204
rect 4016 2150 4018 2202
rect 4198 2150 4200 2202
rect 3954 2148 3960 2150
rect 4016 2148 4040 2150
rect 4096 2148 4120 2150
rect 4176 2148 4200 2150
rect 4256 2148 4262 2150
rect 3954 2139 4262 2148
rect 5517 2204 5825 2213
rect 5517 2202 5523 2204
rect 5579 2202 5603 2204
rect 5659 2202 5683 2204
rect 5739 2202 5763 2204
rect 5819 2202 5825 2204
rect 5579 2150 5581 2202
rect 5761 2150 5763 2202
rect 5517 2148 5523 2150
rect 5579 2148 5603 2150
rect 5659 2148 5683 2150
rect 5739 2148 5763 2150
rect 5819 2148 5825 2150
rect 5517 2139 5825 2148
rect 7080 2204 7388 2213
rect 7080 2202 7086 2204
rect 7142 2202 7166 2204
rect 7222 2202 7246 2204
rect 7302 2202 7326 2204
rect 7382 2202 7388 2204
rect 7142 2150 7144 2202
rect 7324 2150 7326 2202
rect 7080 2148 7086 2150
rect 7142 2148 7166 2150
rect 7222 2148 7246 2150
rect 7302 2148 7326 2150
rect 7382 2148 7388 2150
rect 7080 2139 7388 2148
<< via2 >>
rect 1737 8186 1793 8188
rect 1817 8186 1873 8188
rect 1897 8186 1953 8188
rect 1977 8186 2033 8188
rect 1737 8134 1783 8186
rect 1783 8134 1793 8186
rect 1817 8134 1847 8186
rect 1847 8134 1859 8186
rect 1859 8134 1873 8186
rect 1897 8134 1911 8186
rect 1911 8134 1923 8186
rect 1923 8134 1953 8186
rect 1977 8134 1987 8186
rect 1987 8134 2033 8186
rect 1737 8132 1793 8134
rect 1817 8132 1873 8134
rect 1897 8132 1953 8134
rect 1977 8132 2033 8134
rect 3300 8186 3356 8188
rect 3380 8186 3436 8188
rect 3460 8186 3516 8188
rect 3540 8186 3596 8188
rect 3300 8134 3346 8186
rect 3346 8134 3356 8186
rect 3380 8134 3410 8186
rect 3410 8134 3422 8186
rect 3422 8134 3436 8186
rect 3460 8134 3474 8186
rect 3474 8134 3486 8186
rect 3486 8134 3516 8186
rect 3540 8134 3550 8186
rect 3550 8134 3596 8186
rect 3300 8132 3356 8134
rect 3380 8132 3436 8134
rect 3460 8132 3516 8134
rect 3540 8132 3596 8134
rect 4863 8186 4919 8188
rect 4943 8186 4999 8188
rect 5023 8186 5079 8188
rect 5103 8186 5159 8188
rect 4863 8134 4909 8186
rect 4909 8134 4919 8186
rect 4943 8134 4973 8186
rect 4973 8134 4985 8186
rect 4985 8134 4999 8186
rect 5023 8134 5037 8186
rect 5037 8134 5049 8186
rect 5049 8134 5079 8186
rect 5103 8134 5113 8186
rect 5113 8134 5159 8186
rect 4863 8132 4919 8134
rect 4943 8132 4999 8134
rect 5023 8132 5079 8134
rect 5103 8132 5159 8134
rect 6426 8186 6482 8188
rect 6506 8186 6562 8188
rect 6586 8186 6642 8188
rect 6666 8186 6722 8188
rect 6426 8134 6472 8186
rect 6472 8134 6482 8186
rect 6506 8134 6536 8186
rect 6536 8134 6548 8186
rect 6548 8134 6562 8186
rect 6586 8134 6600 8186
rect 6600 8134 6612 8186
rect 6612 8134 6642 8186
rect 6666 8134 6676 8186
rect 6676 8134 6722 8186
rect 6426 8132 6482 8134
rect 6506 8132 6562 8134
rect 6586 8132 6642 8134
rect 6666 8132 6722 8134
rect 2397 7642 2453 7644
rect 2477 7642 2533 7644
rect 2557 7642 2613 7644
rect 2637 7642 2693 7644
rect 2397 7590 2443 7642
rect 2443 7590 2453 7642
rect 2477 7590 2507 7642
rect 2507 7590 2519 7642
rect 2519 7590 2533 7642
rect 2557 7590 2571 7642
rect 2571 7590 2583 7642
rect 2583 7590 2613 7642
rect 2637 7590 2647 7642
rect 2647 7590 2693 7642
rect 2397 7588 2453 7590
rect 2477 7588 2533 7590
rect 2557 7588 2613 7590
rect 2637 7588 2693 7590
rect 3960 7642 4016 7644
rect 4040 7642 4096 7644
rect 4120 7642 4176 7644
rect 4200 7642 4256 7644
rect 3960 7590 4006 7642
rect 4006 7590 4016 7642
rect 4040 7590 4070 7642
rect 4070 7590 4082 7642
rect 4082 7590 4096 7642
rect 4120 7590 4134 7642
rect 4134 7590 4146 7642
rect 4146 7590 4176 7642
rect 4200 7590 4210 7642
rect 4210 7590 4256 7642
rect 3960 7588 4016 7590
rect 4040 7588 4096 7590
rect 4120 7588 4176 7590
rect 4200 7588 4256 7590
rect 5523 7642 5579 7644
rect 5603 7642 5659 7644
rect 5683 7642 5739 7644
rect 5763 7642 5819 7644
rect 5523 7590 5569 7642
rect 5569 7590 5579 7642
rect 5603 7590 5633 7642
rect 5633 7590 5645 7642
rect 5645 7590 5659 7642
rect 5683 7590 5697 7642
rect 5697 7590 5709 7642
rect 5709 7590 5739 7642
rect 5763 7590 5773 7642
rect 5773 7590 5819 7642
rect 5523 7588 5579 7590
rect 5603 7588 5659 7590
rect 5683 7588 5739 7590
rect 5763 7588 5819 7590
rect 7086 7642 7142 7644
rect 7166 7642 7222 7644
rect 7246 7642 7302 7644
rect 7326 7642 7382 7644
rect 7086 7590 7132 7642
rect 7132 7590 7142 7642
rect 7166 7590 7196 7642
rect 7196 7590 7208 7642
rect 7208 7590 7222 7642
rect 7246 7590 7260 7642
rect 7260 7590 7272 7642
rect 7272 7590 7302 7642
rect 7326 7590 7336 7642
rect 7336 7590 7382 7642
rect 7086 7588 7142 7590
rect 7166 7588 7222 7590
rect 7246 7588 7302 7590
rect 7326 7588 7382 7590
rect 1737 7098 1793 7100
rect 1817 7098 1873 7100
rect 1897 7098 1953 7100
rect 1977 7098 2033 7100
rect 1737 7046 1783 7098
rect 1783 7046 1793 7098
rect 1817 7046 1847 7098
rect 1847 7046 1859 7098
rect 1859 7046 1873 7098
rect 1897 7046 1911 7098
rect 1911 7046 1923 7098
rect 1923 7046 1953 7098
rect 1977 7046 1987 7098
rect 1987 7046 2033 7098
rect 1737 7044 1793 7046
rect 1817 7044 1873 7046
rect 1897 7044 1953 7046
rect 1977 7044 2033 7046
rect 3300 7098 3356 7100
rect 3380 7098 3436 7100
rect 3460 7098 3516 7100
rect 3540 7098 3596 7100
rect 3300 7046 3346 7098
rect 3346 7046 3356 7098
rect 3380 7046 3410 7098
rect 3410 7046 3422 7098
rect 3422 7046 3436 7098
rect 3460 7046 3474 7098
rect 3474 7046 3486 7098
rect 3486 7046 3516 7098
rect 3540 7046 3550 7098
rect 3550 7046 3596 7098
rect 3300 7044 3356 7046
rect 3380 7044 3436 7046
rect 3460 7044 3516 7046
rect 3540 7044 3596 7046
rect 4863 7098 4919 7100
rect 4943 7098 4999 7100
rect 5023 7098 5079 7100
rect 5103 7098 5159 7100
rect 4863 7046 4909 7098
rect 4909 7046 4919 7098
rect 4943 7046 4973 7098
rect 4973 7046 4985 7098
rect 4985 7046 4999 7098
rect 5023 7046 5037 7098
rect 5037 7046 5049 7098
rect 5049 7046 5079 7098
rect 5103 7046 5113 7098
rect 5113 7046 5159 7098
rect 4863 7044 4919 7046
rect 4943 7044 4999 7046
rect 5023 7044 5079 7046
rect 5103 7044 5159 7046
rect 6426 7098 6482 7100
rect 6506 7098 6562 7100
rect 6586 7098 6642 7100
rect 6666 7098 6722 7100
rect 6426 7046 6472 7098
rect 6472 7046 6482 7098
rect 6506 7046 6536 7098
rect 6536 7046 6548 7098
rect 6548 7046 6562 7098
rect 6586 7046 6600 7098
rect 6600 7046 6612 7098
rect 6612 7046 6642 7098
rect 6666 7046 6676 7098
rect 6676 7046 6722 7098
rect 6426 7044 6482 7046
rect 6506 7044 6562 7046
rect 6586 7044 6642 7046
rect 6666 7044 6722 7046
rect 2397 6554 2453 6556
rect 2477 6554 2533 6556
rect 2557 6554 2613 6556
rect 2637 6554 2693 6556
rect 2397 6502 2443 6554
rect 2443 6502 2453 6554
rect 2477 6502 2507 6554
rect 2507 6502 2519 6554
rect 2519 6502 2533 6554
rect 2557 6502 2571 6554
rect 2571 6502 2583 6554
rect 2583 6502 2613 6554
rect 2637 6502 2647 6554
rect 2647 6502 2693 6554
rect 2397 6500 2453 6502
rect 2477 6500 2533 6502
rect 2557 6500 2613 6502
rect 2637 6500 2693 6502
rect 3960 6554 4016 6556
rect 4040 6554 4096 6556
rect 4120 6554 4176 6556
rect 4200 6554 4256 6556
rect 3960 6502 4006 6554
rect 4006 6502 4016 6554
rect 4040 6502 4070 6554
rect 4070 6502 4082 6554
rect 4082 6502 4096 6554
rect 4120 6502 4134 6554
rect 4134 6502 4146 6554
rect 4146 6502 4176 6554
rect 4200 6502 4210 6554
rect 4210 6502 4256 6554
rect 3960 6500 4016 6502
rect 4040 6500 4096 6502
rect 4120 6500 4176 6502
rect 4200 6500 4256 6502
rect 5523 6554 5579 6556
rect 5603 6554 5659 6556
rect 5683 6554 5739 6556
rect 5763 6554 5819 6556
rect 5523 6502 5569 6554
rect 5569 6502 5579 6554
rect 5603 6502 5633 6554
rect 5633 6502 5645 6554
rect 5645 6502 5659 6554
rect 5683 6502 5697 6554
rect 5697 6502 5709 6554
rect 5709 6502 5739 6554
rect 5763 6502 5773 6554
rect 5773 6502 5819 6554
rect 5523 6500 5579 6502
rect 5603 6500 5659 6502
rect 5683 6500 5739 6502
rect 5763 6500 5819 6502
rect 7086 6554 7142 6556
rect 7166 6554 7222 6556
rect 7246 6554 7302 6556
rect 7326 6554 7382 6556
rect 7086 6502 7132 6554
rect 7132 6502 7142 6554
rect 7166 6502 7196 6554
rect 7196 6502 7208 6554
rect 7208 6502 7222 6554
rect 7246 6502 7260 6554
rect 7260 6502 7272 6554
rect 7272 6502 7302 6554
rect 7326 6502 7336 6554
rect 7336 6502 7382 6554
rect 7086 6500 7142 6502
rect 7166 6500 7222 6502
rect 7246 6500 7302 6502
rect 7326 6500 7382 6502
rect 1737 6010 1793 6012
rect 1817 6010 1873 6012
rect 1897 6010 1953 6012
rect 1977 6010 2033 6012
rect 1737 5958 1783 6010
rect 1783 5958 1793 6010
rect 1817 5958 1847 6010
rect 1847 5958 1859 6010
rect 1859 5958 1873 6010
rect 1897 5958 1911 6010
rect 1911 5958 1923 6010
rect 1923 5958 1953 6010
rect 1977 5958 1987 6010
rect 1987 5958 2033 6010
rect 1737 5956 1793 5958
rect 1817 5956 1873 5958
rect 1897 5956 1953 5958
rect 1977 5956 2033 5958
rect 3300 6010 3356 6012
rect 3380 6010 3436 6012
rect 3460 6010 3516 6012
rect 3540 6010 3596 6012
rect 3300 5958 3346 6010
rect 3346 5958 3356 6010
rect 3380 5958 3410 6010
rect 3410 5958 3422 6010
rect 3422 5958 3436 6010
rect 3460 5958 3474 6010
rect 3474 5958 3486 6010
rect 3486 5958 3516 6010
rect 3540 5958 3550 6010
rect 3550 5958 3596 6010
rect 3300 5956 3356 5958
rect 3380 5956 3436 5958
rect 3460 5956 3516 5958
rect 3540 5956 3596 5958
rect 4863 6010 4919 6012
rect 4943 6010 4999 6012
rect 5023 6010 5079 6012
rect 5103 6010 5159 6012
rect 4863 5958 4909 6010
rect 4909 5958 4919 6010
rect 4943 5958 4973 6010
rect 4973 5958 4985 6010
rect 4985 5958 4999 6010
rect 5023 5958 5037 6010
rect 5037 5958 5049 6010
rect 5049 5958 5079 6010
rect 5103 5958 5113 6010
rect 5113 5958 5159 6010
rect 4863 5956 4919 5958
rect 4943 5956 4999 5958
rect 5023 5956 5079 5958
rect 5103 5956 5159 5958
rect 6426 6010 6482 6012
rect 6506 6010 6562 6012
rect 6586 6010 6642 6012
rect 6666 6010 6722 6012
rect 6426 5958 6472 6010
rect 6472 5958 6482 6010
rect 6506 5958 6536 6010
rect 6536 5958 6548 6010
rect 6548 5958 6562 6010
rect 6586 5958 6600 6010
rect 6600 5958 6612 6010
rect 6612 5958 6642 6010
rect 6666 5958 6676 6010
rect 6676 5958 6722 6010
rect 6426 5956 6482 5958
rect 6506 5956 6562 5958
rect 6586 5956 6642 5958
rect 6666 5956 6722 5958
rect 1398 5480 1454 5536
rect 2397 5466 2453 5468
rect 2477 5466 2533 5468
rect 2557 5466 2613 5468
rect 2637 5466 2693 5468
rect 2397 5414 2443 5466
rect 2443 5414 2453 5466
rect 2477 5414 2507 5466
rect 2507 5414 2519 5466
rect 2519 5414 2533 5466
rect 2557 5414 2571 5466
rect 2571 5414 2583 5466
rect 2583 5414 2613 5466
rect 2637 5414 2647 5466
rect 2647 5414 2693 5466
rect 2397 5412 2453 5414
rect 2477 5412 2533 5414
rect 2557 5412 2613 5414
rect 2637 5412 2693 5414
rect 846 4972 848 4992
rect 848 4972 900 4992
rect 900 4972 902 4992
rect 846 4936 902 4972
rect 1737 4922 1793 4924
rect 1817 4922 1873 4924
rect 1897 4922 1953 4924
rect 1977 4922 2033 4924
rect 1737 4870 1783 4922
rect 1783 4870 1793 4922
rect 1817 4870 1847 4922
rect 1847 4870 1859 4922
rect 1859 4870 1873 4922
rect 1897 4870 1911 4922
rect 1911 4870 1923 4922
rect 1923 4870 1953 4922
rect 1977 4870 1987 4922
rect 1987 4870 2033 4922
rect 1737 4868 1793 4870
rect 1817 4868 1873 4870
rect 1897 4868 1953 4870
rect 1977 4868 2033 4870
rect 3960 5466 4016 5468
rect 4040 5466 4096 5468
rect 4120 5466 4176 5468
rect 4200 5466 4256 5468
rect 3960 5414 4006 5466
rect 4006 5414 4016 5466
rect 4040 5414 4070 5466
rect 4070 5414 4082 5466
rect 4082 5414 4096 5466
rect 4120 5414 4134 5466
rect 4134 5414 4146 5466
rect 4146 5414 4176 5466
rect 4200 5414 4210 5466
rect 4210 5414 4256 5466
rect 3960 5412 4016 5414
rect 4040 5412 4096 5414
rect 4120 5412 4176 5414
rect 4200 5412 4256 5414
rect 5523 5466 5579 5468
rect 5603 5466 5659 5468
rect 5683 5466 5739 5468
rect 5763 5466 5819 5468
rect 5523 5414 5569 5466
rect 5569 5414 5579 5466
rect 5603 5414 5633 5466
rect 5633 5414 5645 5466
rect 5645 5414 5659 5466
rect 5683 5414 5697 5466
rect 5697 5414 5709 5466
rect 5709 5414 5739 5466
rect 5763 5414 5773 5466
rect 5773 5414 5819 5466
rect 5523 5412 5579 5414
rect 5603 5412 5659 5414
rect 5683 5412 5739 5414
rect 5763 5412 5819 5414
rect 7470 5516 7472 5536
rect 7472 5516 7524 5536
rect 7524 5516 7526 5536
rect 7470 5480 7526 5516
rect 7086 5466 7142 5468
rect 7166 5466 7222 5468
rect 7246 5466 7302 5468
rect 7326 5466 7382 5468
rect 7086 5414 7132 5466
rect 7132 5414 7142 5466
rect 7166 5414 7196 5466
rect 7196 5414 7208 5466
rect 7208 5414 7222 5466
rect 7246 5414 7260 5466
rect 7260 5414 7272 5466
rect 7272 5414 7302 5466
rect 7326 5414 7336 5466
rect 7336 5414 7382 5466
rect 7086 5412 7142 5414
rect 7166 5412 7222 5414
rect 7246 5412 7302 5414
rect 7326 5412 7382 5414
rect 3300 4922 3356 4924
rect 3380 4922 3436 4924
rect 3460 4922 3516 4924
rect 3540 4922 3596 4924
rect 3300 4870 3346 4922
rect 3346 4870 3356 4922
rect 3380 4870 3410 4922
rect 3410 4870 3422 4922
rect 3422 4870 3436 4922
rect 3460 4870 3474 4922
rect 3474 4870 3486 4922
rect 3486 4870 3516 4922
rect 3540 4870 3550 4922
rect 3550 4870 3596 4922
rect 3300 4868 3356 4870
rect 3380 4868 3436 4870
rect 3460 4868 3516 4870
rect 3540 4868 3596 4870
rect 4863 4922 4919 4924
rect 4943 4922 4999 4924
rect 5023 4922 5079 4924
rect 5103 4922 5159 4924
rect 4863 4870 4909 4922
rect 4909 4870 4919 4922
rect 4943 4870 4973 4922
rect 4973 4870 4985 4922
rect 4985 4870 4999 4922
rect 5023 4870 5037 4922
rect 5037 4870 5049 4922
rect 5049 4870 5079 4922
rect 5103 4870 5113 4922
rect 5113 4870 5159 4922
rect 4863 4868 4919 4870
rect 4943 4868 4999 4870
rect 5023 4868 5079 4870
rect 5103 4868 5159 4870
rect 6426 4922 6482 4924
rect 6506 4922 6562 4924
rect 6586 4922 6642 4924
rect 6666 4922 6722 4924
rect 6426 4870 6472 4922
rect 6472 4870 6482 4922
rect 6506 4870 6536 4922
rect 6536 4870 6548 4922
rect 6548 4870 6562 4922
rect 6586 4870 6600 4922
rect 6600 4870 6612 4922
rect 6612 4870 6642 4922
rect 6666 4870 6676 4922
rect 6676 4870 6722 4922
rect 6426 4868 6482 4870
rect 6506 4868 6562 4870
rect 6586 4868 6642 4870
rect 6666 4868 6722 4870
rect 7010 4800 7066 4856
rect 2397 4378 2453 4380
rect 2477 4378 2533 4380
rect 2557 4378 2613 4380
rect 2637 4378 2693 4380
rect 2397 4326 2443 4378
rect 2443 4326 2453 4378
rect 2477 4326 2507 4378
rect 2507 4326 2519 4378
rect 2519 4326 2533 4378
rect 2557 4326 2571 4378
rect 2571 4326 2583 4378
rect 2583 4326 2613 4378
rect 2637 4326 2647 4378
rect 2647 4326 2693 4378
rect 2397 4324 2453 4326
rect 2477 4324 2533 4326
rect 2557 4324 2613 4326
rect 2637 4324 2693 4326
rect 3960 4378 4016 4380
rect 4040 4378 4096 4380
rect 4120 4378 4176 4380
rect 4200 4378 4256 4380
rect 3960 4326 4006 4378
rect 4006 4326 4016 4378
rect 4040 4326 4070 4378
rect 4070 4326 4082 4378
rect 4082 4326 4096 4378
rect 4120 4326 4134 4378
rect 4134 4326 4146 4378
rect 4146 4326 4176 4378
rect 4200 4326 4210 4378
rect 4210 4326 4256 4378
rect 3960 4324 4016 4326
rect 4040 4324 4096 4326
rect 4120 4324 4176 4326
rect 4200 4324 4256 4326
rect 5523 4378 5579 4380
rect 5603 4378 5659 4380
rect 5683 4378 5739 4380
rect 5763 4378 5819 4380
rect 5523 4326 5569 4378
rect 5569 4326 5579 4378
rect 5603 4326 5633 4378
rect 5633 4326 5645 4378
rect 5645 4326 5659 4378
rect 5683 4326 5697 4378
rect 5697 4326 5709 4378
rect 5709 4326 5739 4378
rect 5763 4326 5773 4378
rect 5773 4326 5819 4378
rect 5523 4324 5579 4326
rect 5603 4324 5659 4326
rect 5683 4324 5739 4326
rect 5763 4324 5819 4326
rect 7086 4378 7142 4380
rect 7166 4378 7222 4380
rect 7246 4378 7302 4380
rect 7326 4378 7382 4380
rect 7086 4326 7132 4378
rect 7132 4326 7142 4378
rect 7166 4326 7196 4378
rect 7196 4326 7208 4378
rect 7208 4326 7222 4378
rect 7246 4326 7260 4378
rect 7260 4326 7272 4378
rect 7272 4326 7302 4378
rect 7326 4326 7336 4378
rect 7336 4326 7382 4378
rect 7086 4324 7142 4326
rect 7166 4324 7222 4326
rect 7246 4324 7302 4326
rect 7326 4324 7382 4326
rect 846 4256 902 4312
rect 1737 3834 1793 3836
rect 1817 3834 1873 3836
rect 1897 3834 1953 3836
rect 1977 3834 2033 3836
rect 1737 3782 1783 3834
rect 1783 3782 1793 3834
rect 1817 3782 1847 3834
rect 1847 3782 1859 3834
rect 1859 3782 1873 3834
rect 1897 3782 1911 3834
rect 1911 3782 1923 3834
rect 1923 3782 1953 3834
rect 1977 3782 1987 3834
rect 1987 3782 2033 3834
rect 1737 3780 1793 3782
rect 1817 3780 1873 3782
rect 1897 3780 1953 3782
rect 1977 3780 2033 3782
rect 3300 3834 3356 3836
rect 3380 3834 3436 3836
rect 3460 3834 3516 3836
rect 3540 3834 3596 3836
rect 3300 3782 3346 3834
rect 3346 3782 3356 3834
rect 3380 3782 3410 3834
rect 3410 3782 3422 3834
rect 3422 3782 3436 3834
rect 3460 3782 3474 3834
rect 3474 3782 3486 3834
rect 3486 3782 3516 3834
rect 3540 3782 3550 3834
rect 3550 3782 3596 3834
rect 3300 3780 3356 3782
rect 3380 3780 3436 3782
rect 3460 3780 3516 3782
rect 3540 3780 3596 3782
rect 4863 3834 4919 3836
rect 4943 3834 4999 3836
rect 5023 3834 5079 3836
rect 5103 3834 5159 3836
rect 4863 3782 4909 3834
rect 4909 3782 4919 3834
rect 4943 3782 4973 3834
rect 4973 3782 4985 3834
rect 4985 3782 4999 3834
rect 5023 3782 5037 3834
rect 5037 3782 5049 3834
rect 5049 3782 5079 3834
rect 5103 3782 5113 3834
rect 5113 3782 5159 3834
rect 4863 3780 4919 3782
rect 4943 3780 4999 3782
rect 5023 3780 5079 3782
rect 5103 3780 5159 3782
rect 6426 3834 6482 3836
rect 6506 3834 6562 3836
rect 6586 3834 6642 3836
rect 6666 3834 6722 3836
rect 6426 3782 6472 3834
rect 6472 3782 6482 3834
rect 6506 3782 6536 3834
rect 6536 3782 6548 3834
rect 6548 3782 6562 3834
rect 6586 3782 6600 3834
rect 6600 3782 6612 3834
rect 6612 3782 6642 3834
rect 6666 3782 6676 3834
rect 6676 3782 6722 3834
rect 6426 3780 6482 3782
rect 6506 3780 6562 3782
rect 6586 3780 6642 3782
rect 6666 3780 6722 3782
rect 2397 3290 2453 3292
rect 2477 3290 2533 3292
rect 2557 3290 2613 3292
rect 2637 3290 2693 3292
rect 2397 3238 2443 3290
rect 2443 3238 2453 3290
rect 2477 3238 2507 3290
rect 2507 3238 2519 3290
rect 2519 3238 2533 3290
rect 2557 3238 2571 3290
rect 2571 3238 2583 3290
rect 2583 3238 2613 3290
rect 2637 3238 2647 3290
rect 2647 3238 2693 3290
rect 2397 3236 2453 3238
rect 2477 3236 2533 3238
rect 2557 3236 2613 3238
rect 2637 3236 2693 3238
rect 3960 3290 4016 3292
rect 4040 3290 4096 3292
rect 4120 3290 4176 3292
rect 4200 3290 4256 3292
rect 3960 3238 4006 3290
rect 4006 3238 4016 3290
rect 4040 3238 4070 3290
rect 4070 3238 4082 3290
rect 4082 3238 4096 3290
rect 4120 3238 4134 3290
rect 4134 3238 4146 3290
rect 4146 3238 4176 3290
rect 4200 3238 4210 3290
rect 4210 3238 4256 3290
rect 3960 3236 4016 3238
rect 4040 3236 4096 3238
rect 4120 3236 4176 3238
rect 4200 3236 4256 3238
rect 5523 3290 5579 3292
rect 5603 3290 5659 3292
rect 5683 3290 5739 3292
rect 5763 3290 5819 3292
rect 5523 3238 5569 3290
rect 5569 3238 5579 3290
rect 5603 3238 5633 3290
rect 5633 3238 5645 3290
rect 5645 3238 5659 3290
rect 5683 3238 5697 3290
rect 5697 3238 5709 3290
rect 5709 3238 5739 3290
rect 5763 3238 5773 3290
rect 5773 3238 5819 3290
rect 5523 3236 5579 3238
rect 5603 3236 5659 3238
rect 5683 3236 5739 3238
rect 5763 3236 5819 3238
rect 7086 3290 7142 3292
rect 7166 3290 7222 3292
rect 7246 3290 7302 3292
rect 7326 3290 7382 3292
rect 7086 3238 7132 3290
rect 7132 3238 7142 3290
rect 7166 3238 7196 3290
rect 7196 3238 7208 3290
rect 7208 3238 7222 3290
rect 7246 3238 7260 3290
rect 7260 3238 7272 3290
rect 7272 3238 7302 3290
rect 7326 3238 7336 3290
rect 7336 3238 7382 3290
rect 7086 3236 7142 3238
rect 7166 3236 7222 3238
rect 7246 3236 7302 3238
rect 7326 3236 7382 3238
rect 1737 2746 1793 2748
rect 1817 2746 1873 2748
rect 1897 2746 1953 2748
rect 1977 2746 2033 2748
rect 1737 2694 1783 2746
rect 1783 2694 1793 2746
rect 1817 2694 1847 2746
rect 1847 2694 1859 2746
rect 1859 2694 1873 2746
rect 1897 2694 1911 2746
rect 1911 2694 1923 2746
rect 1923 2694 1953 2746
rect 1977 2694 1987 2746
rect 1987 2694 2033 2746
rect 1737 2692 1793 2694
rect 1817 2692 1873 2694
rect 1897 2692 1953 2694
rect 1977 2692 2033 2694
rect 3300 2746 3356 2748
rect 3380 2746 3436 2748
rect 3460 2746 3516 2748
rect 3540 2746 3596 2748
rect 3300 2694 3346 2746
rect 3346 2694 3356 2746
rect 3380 2694 3410 2746
rect 3410 2694 3422 2746
rect 3422 2694 3436 2746
rect 3460 2694 3474 2746
rect 3474 2694 3486 2746
rect 3486 2694 3516 2746
rect 3540 2694 3550 2746
rect 3550 2694 3596 2746
rect 3300 2692 3356 2694
rect 3380 2692 3436 2694
rect 3460 2692 3516 2694
rect 3540 2692 3596 2694
rect 4863 2746 4919 2748
rect 4943 2746 4999 2748
rect 5023 2746 5079 2748
rect 5103 2746 5159 2748
rect 4863 2694 4909 2746
rect 4909 2694 4919 2746
rect 4943 2694 4973 2746
rect 4973 2694 4985 2746
rect 4985 2694 4999 2746
rect 5023 2694 5037 2746
rect 5037 2694 5049 2746
rect 5049 2694 5079 2746
rect 5103 2694 5113 2746
rect 5113 2694 5159 2746
rect 4863 2692 4919 2694
rect 4943 2692 4999 2694
rect 5023 2692 5079 2694
rect 5103 2692 5159 2694
rect 6426 2746 6482 2748
rect 6506 2746 6562 2748
rect 6586 2746 6642 2748
rect 6666 2746 6722 2748
rect 6426 2694 6472 2746
rect 6472 2694 6482 2746
rect 6506 2694 6536 2746
rect 6536 2694 6548 2746
rect 6548 2694 6562 2746
rect 6586 2694 6600 2746
rect 6600 2694 6612 2746
rect 6612 2694 6642 2746
rect 6666 2694 6676 2746
rect 6676 2694 6722 2746
rect 6426 2692 6482 2694
rect 6506 2692 6562 2694
rect 6586 2692 6642 2694
rect 6666 2692 6722 2694
rect 2397 2202 2453 2204
rect 2477 2202 2533 2204
rect 2557 2202 2613 2204
rect 2637 2202 2693 2204
rect 2397 2150 2443 2202
rect 2443 2150 2453 2202
rect 2477 2150 2507 2202
rect 2507 2150 2519 2202
rect 2519 2150 2533 2202
rect 2557 2150 2571 2202
rect 2571 2150 2583 2202
rect 2583 2150 2613 2202
rect 2637 2150 2647 2202
rect 2647 2150 2693 2202
rect 2397 2148 2453 2150
rect 2477 2148 2533 2150
rect 2557 2148 2613 2150
rect 2637 2148 2693 2150
rect 3960 2202 4016 2204
rect 4040 2202 4096 2204
rect 4120 2202 4176 2204
rect 4200 2202 4256 2204
rect 3960 2150 4006 2202
rect 4006 2150 4016 2202
rect 4040 2150 4070 2202
rect 4070 2150 4082 2202
rect 4082 2150 4096 2202
rect 4120 2150 4134 2202
rect 4134 2150 4146 2202
rect 4146 2150 4176 2202
rect 4200 2150 4210 2202
rect 4210 2150 4256 2202
rect 3960 2148 4016 2150
rect 4040 2148 4096 2150
rect 4120 2148 4176 2150
rect 4200 2148 4256 2150
rect 5523 2202 5579 2204
rect 5603 2202 5659 2204
rect 5683 2202 5739 2204
rect 5763 2202 5819 2204
rect 5523 2150 5569 2202
rect 5569 2150 5579 2202
rect 5603 2150 5633 2202
rect 5633 2150 5645 2202
rect 5645 2150 5659 2202
rect 5683 2150 5697 2202
rect 5697 2150 5709 2202
rect 5709 2150 5739 2202
rect 5763 2150 5773 2202
rect 5773 2150 5819 2202
rect 5523 2148 5579 2150
rect 5603 2148 5659 2150
rect 5683 2148 5739 2150
rect 5763 2148 5819 2150
rect 7086 2202 7142 2204
rect 7166 2202 7222 2204
rect 7246 2202 7302 2204
rect 7326 2202 7382 2204
rect 7086 2150 7132 2202
rect 7132 2150 7142 2202
rect 7166 2150 7196 2202
rect 7196 2150 7208 2202
rect 7208 2150 7222 2202
rect 7246 2150 7260 2202
rect 7260 2150 7272 2202
rect 7272 2150 7302 2202
rect 7326 2150 7336 2202
rect 7336 2150 7382 2202
rect 7086 2148 7142 2150
rect 7166 2148 7222 2150
rect 7246 2148 7302 2150
rect 7326 2148 7382 2150
<< metal3 >>
rect 1727 8192 2043 8193
rect 1727 8128 1733 8192
rect 1797 8128 1813 8192
rect 1877 8128 1893 8192
rect 1957 8128 1973 8192
rect 2037 8128 2043 8192
rect 1727 8127 2043 8128
rect 3290 8192 3606 8193
rect 3290 8128 3296 8192
rect 3360 8128 3376 8192
rect 3440 8128 3456 8192
rect 3520 8128 3536 8192
rect 3600 8128 3606 8192
rect 3290 8127 3606 8128
rect 4853 8192 5169 8193
rect 4853 8128 4859 8192
rect 4923 8128 4939 8192
rect 5003 8128 5019 8192
rect 5083 8128 5099 8192
rect 5163 8128 5169 8192
rect 4853 8127 5169 8128
rect 6416 8192 6732 8193
rect 6416 8128 6422 8192
rect 6486 8128 6502 8192
rect 6566 8128 6582 8192
rect 6646 8128 6662 8192
rect 6726 8128 6732 8192
rect 6416 8127 6732 8128
rect 2387 7648 2703 7649
rect 2387 7584 2393 7648
rect 2457 7584 2473 7648
rect 2537 7584 2553 7648
rect 2617 7584 2633 7648
rect 2697 7584 2703 7648
rect 2387 7583 2703 7584
rect 3950 7648 4266 7649
rect 3950 7584 3956 7648
rect 4020 7584 4036 7648
rect 4100 7584 4116 7648
rect 4180 7584 4196 7648
rect 4260 7584 4266 7648
rect 3950 7583 4266 7584
rect 5513 7648 5829 7649
rect 5513 7584 5519 7648
rect 5583 7584 5599 7648
rect 5663 7584 5679 7648
rect 5743 7584 5759 7648
rect 5823 7584 5829 7648
rect 5513 7583 5829 7584
rect 7076 7648 7392 7649
rect 7076 7584 7082 7648
rect 7146 7584 7162 7648
rect 7226 7584 7242 7648
rect 7306 7584 7322 7648
rect 7386 7584 7392 7648
rect 7076 7583 7392 7584
rect 1727 7104 2043 7105
rect 1727 7040 1733 7104
rect 1797 7040 1813 7104
rect 1877 7040 1893 7104
rect 1957 7040 1973 7104
rect 2037 7040 2043 7104
rect 1727 7039 2043 7040
rect 3290 7104 3606 7105
rect 3290 7040 3296 7104
rect 3360 7040 3376 7104
rect 3440 7040 3456 7104
rect 3520 7040 3536 7104
rect 3600 7040 3606 7104
rect 3290 7039 3606 7040
rect 4853 7104 5169 7105
rect 4853 7040 4859 7104
rect 4923 7040 4939 7104
rect 5003 7040 5019 7104
rect 5083 7040 5099 7104
rect 5163 7040 5169 7104
rect 4853 7039 5169 7040
rect 6416 7104 6732 7105
rect 6416 7040 6422 7104
rect 6486 7040 6502 7104
rect 6566 7040 6582 7104
rect 6646 7040 6662 7104
rect 6726 7040 6732 7104
rect 6416 7039 6732 7040
rect 2387 6560 2703 6561
rect 2387 6496 2393 6560
rect 2457 6496 2473 6560
rect 2537 6496 2553 6560
rect 2617 6496 2633 6560
rect 2697 6496 2703 6560
rect 2387 6495 2703 6496
rect 3950 6560 4266 6561
rect 3950 6496 3956 6560
rect 4020 6496 4036 6560
rect 4100 6496 4116 6560
rect 4180 6496 4196 6560
rect 4260 6496 4266 6560
rect 3950 6495 4266 6496
rect 5513 6560 5829 6561
rect 5513 6496 5519 6560
rect 5583 6496 5599 6560
rect 5663 6496 5679 6560
rect 5743 6496 5759 6560
rect 5823 6496 5829 6560
rect 5513 6495 5829 6496
rect 7076 6560 7392 6561
rect 7076 6496 7082 6560
rect 7146 6496 7162 6560
rect 7226 6496 7242 6560
rect 7306 6496 7322 6560
rect 7386 6496 7392 6560
rect 7076 6495 7392 6496
rect 1727 6016 2043 6017
rect 1727 5952 1733 6016
rect 1797 5952 1813 6016
rect 1877 5952 1893 6016
rect 1957 5952 1973 6016
rect 2037 5952 2043 6016
rect 1727 5951 2043 5952
rect 3290 6016 3606 6017
rect 3290 5952 3296 6016
rect 3360 5952 3376 6016
rect 3440 5952 3456 6016
rect 3520 5952 3536 6016
rect 3600 5952 3606 6016
rect 3290 5951 3606 5952
rect 4853 6016 5169 6017
rect 4853 5952 4859 6016
rect 4923 5952 4939 6016
rect 5003 5952 5019 6016
rect 5083 5952 5099 6016
rect 5163 5952 5169 6016
rect 4853 5951 5169 5952
rect 6416 6016 6732 6017
rect 6416 5952 6422 6016
rect 6486 5952 6502 6016
rect 6566 5952 6582 6016
rect 6646 5952 6662 6016
rect 6726 5952 6732 6016
rect 6416 5951 6732 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 7465 5538 7531 5541
rect 7735 5538 8535 5568
rect 7465 5536 8535 5538
rect 7465 5480 7470 5536
rect 7526 5480 8535 5536
rect 7465 5478 8535 5480
rect 7465 5475 7531 5478
rect 2387 5472 2703 5473
rect 2387 5408 2393 5472
rect 2457 5408 2473 5472
rect 2537 5408 2553 5472
rect 2617 5408 2633 5472
rect 2697 5408 2703 5472
rect 2387 5407 2703 5408
rect 3950 5472 4266 5473
rect 3950 5408 3956 5472
rect 4020 5408 4036 5472
rect 4100 5408 4116 5472
rect 4180 5408 4196 5472
rect 4260 5408 4266 5472
rect 3950 5407 4266 5408
rect 5513 5472 5829 5473
rect 5513 5408 5519 5472
rect 5583 5408 5599 5472
rect 5663 5408 5679 5472
rect 5743 5408 5759 5472
rect 5823 5408 5829 5472
rect 5513 5407 5829 5408
rect 7076 5472 7392 5473
rect 7076 5408 7082 5472
rect 7146 5408 7162 5472
rect 7226 5408 7242 5472
rect 7306 5408 7322 5472
rect 7386 5408 7392 5472
rect 7735 5448 8535 5478
rect 7076 5407 7392 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 1727 4928 2043 4929
rect 1727 4864 1733 4928
rect 1797 4864 1813 4928
rect 1877 4864 1893 4928
rect 1957 4864 1973 4928
rect 2037 4864 2043 4928
rect 1727 4863 2043 4864
rect 3290 4928 3606 4929
rect 3290 4864 3296 4928
rect 3360 4864 3376 4928
rect 3440 4864 3456 4928
rect 3520 4864 3536 4928
rect 3600 4864 3606 4928
rect 3290 4863 3606 4864
rect 4853 4928 5169 4929
rect 4853 4864 4859 4928
rect 4923 4864 4939 4928
rect 5003 4864 5019 4928
rect 5083 4864 5099 4928
rect 5163 4864 5169 4928
rect 4853 4863 5169 4864
rect 6416 4928 6732 4929
rect 6416 4864 6422 4928
rect 6486 4864 6502 4928
rect 6566 4864 6582 4928
rect 6646 4864 6662 4928
rect 6726 4864 6732 4928
rect 6416 4863 6732 4864
rect 7005 4858 7071 4861
rect 7735 4858 8535 4888
rect 7005 4856 8535 4858
rect 7005 4800 7010 4856
rect 7066 4800 8535 4856
rect 7005 4798 8535 4800
rect 0 4768 800 4798
rect 7005 4795 7071 4798
rect 7735 4768 8535 4798
rect 2387 4384 2703 4385
rect 2387 4320 2393 4384
rect 2457 4320 2473 4384
rect 2537 4320 2553 4384
rect 2617 4320 2633 4384
rect 2697 4320 2703 4384
rect 2387 4319 2703 4320
rect 3950 4384 4266 4385
rect 3950 4320 3956 4384
rect 4020 4320 4036 4384
rect 4100 4320 4116 4384
rect 4180 4320 4196 4384
rect 4260 4320 4266 4384
rect 3950 4319 4266 4320
rect 5513 4384 5829 4385
rect 5513 4320 5519 4384
rect 5583 4320 5599 4384
rect 5663 4320 5679 4384
rect 5743 4320 5759 4384
rect 5823 4320 5829 4384
rect 5513 4319 5829 4320
rect 7076 4384 7392 4385
rect 7076 4320 7082 4384
rect 7146 4320 7162 4384
rect 7226 4320 7242 4384
rect 7306 4320 7322 4384
rect 7386 4320 7392 4384
rect 7076 4319 7392 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 0 4088 800 4118
rect 1727 3840 2043 3841
rect 1727 3776 1733 3840
rect 1797 3776 1813 3840
rect 1877 3776 1893 3840
rect 1957 3776 1973 3840
rect 2037 3776 2043 3840
rect 1727 3775 2043 3776
rect 3290 3840 3606 3841
rect 3290 3776 3296 3840
rect 3360 3776 3376 3840
rect 3440 3776 3456 3840
rect 3520 3776 3536 3840
rect 3600 3776 3606 3840
rect 3290 3775 3606 3776
rect 4853 3840 5169 3841
rect 4853 3776 4859 3840
rect 4923 3776 4939 3840
rect 5003 3776 5019 3840
rect 5083 3776 5099 3840
rect 5163 3776 5169 3840
rect 4853 3775 5169 3776
rect 6416 3840 6732 3841
rect 6416 3776 6422 3840
rect 6486 3776 6502 3840
rect 6566 3776 6582 3840
rect 6646 3776 6662 3840
rect 6726 3776 6732 3840
rect 6416 3775 6732 3776
rect 2387 3296 2703 3297
rect 2387 3232 2393 3296
rect 2457 3232 2473 3296
rect 2537 3232 2553 3296
rect 2617 3232 2633 3296
rect 2697 3232 2703 3296
rect 2387 3231 2703 3232
rect 3950 3296 4266 3297
rect 3950 3232 3956 3296
rect 4020 3232 4036 3296
rect 4100 3232 4116 3296
rect 4180 3232 4196 3296
rect 4260 3232 4266 3296
rect 3950 3231 4266 3232
rect 5513 3296 5829 3297
rect 5513 3232 5519 3296
rect 5583 3232 5599 3296
rect 5663 3232 5679 3296
rect 5743 3232 5759 3296
rect 5823 3232 5829 3296
rect 5513 3231 5829 3232
rect 7076 3296 7392 3297
rect 7076 3232 7082 3296
rect 7146 3232 7162 3296
rect 7226 3232 7242 3296
rect 7306 3232 7322 3296
rect 7386 3232 7392 3296
rect 7076 3231 7392 3232
rect 1727 2752 2043 2753
rect 1727 2688 1733 2752
rect 1797 2688 1813 2752
rect 1877 2688 1893 2752
rect 1957 2688 1973 2752
rect 2037 2688 2043 2752
rect 1727 2687 2043 2688
rect 3290 2752 3606 2753
rect 3290 2688 3296 2752
rect 3360 2688 3376 2752
rect 3440 2688 3456 2752
rect 3520 2688 3536 2752
rect 3600 2688 3606 2752
rect 3290 2687 3606 2688
rect 4853 2752 5169 2753
rect 4853 2688 4859 2752
rect 4923 2688 4939 2752
rect 5003 2688 5019 2752
rect 5083 2688 5099 2752
rect 5163 2688 5169 2752
rect 4853 2687 5169 2688
rect 6416 2752 6732 2753
rect 6416 2688 6422 2752
rect 6486 2688 6502 2752
rect 6566 2688 6582 2752
rect 6646 2688 6662 2752
rect 6726 2688 6732 2752
rect 6416 2687 6732 2688
rect 2387 2208 2703 2209
rect 2387 2144 2393 2208
rect 2457 2144 2473 2208
rect 2537 2144 2553 2208
rect 2617 2144 2633 2208
rect 2697 2144 2703 2208
rect 2387 2143 2703 2144
rect 3950 2208 4266 2209
rect 3950 2144 3956 2208
rect 4020 2144 4036 2208
rect 4100 2144 4116 2208
rect 4180 2144 4196 2208
rect 4260 2144 4266 2208
rect 3950 2143 4266 2144
rect 5513 2208 5829 2209
rect 5513 2144 5519 2208
rect 5583 2144 5599 2208
rect 5663 2144 5679 2208
rect 5743 2144 5759 2208
rect 5823 2144 5829 2208
rect 5513 2143 5829 2144
rect 7076 2208 7392 2209
rect 7076 2144 7082 2208
rect 7146 2144 7162 2208
rect 7226 2144 7242 2208
rect 7306 2144 7322 2208
rect 7386 2144 7392 2208
rect 7076 2143 7392 2144
<< via3 >>
rect 1733 8188 1797 8192
rect 1733 8132 1737 8188
rect 1737 8132 1793 8188
rect 1793 8132 1797 8188
rect 1733 8128 1797 8132
rect 1813 8188 1877 8192
rect 1813 8132 1817 8188
rect 1817 8132 1873 8188
rect 1873 8132 1877 8188
rect 1813 8128 1877 8132
rect 1893 8188 1957 8192
rect 1893 8132 1897 8188
rect 1897 8132 1953 8188
rect 1953 8132 1957 8188
rect 1893 8128 1957 8132
rect 1973 8188 2037 8192
rect 1973 8132 1977 8188
rect 1977 8132 2033 8188
rect 2033 8132 2037 8188
rect 1973 8128 2037 8132
rect 3296 8188 3360 8192
rect 3296 8132 3300 8188
rect 3300 8132 3356 8188
rect 3356 8132 3360 8188
rect 3296 8128 3360 8132
rect 3376 8188 3440 8192
rect 3376 8132 3380 8188
rect 3380 8132 3436 8188
rect 3436 8132 3440 8188
rect 3376 8128 3440 8132
rect 3456 8188 3520 8192
rect 3456 8132 3460 8188
rect 3460 8132 3516 8188
rect 3516 8132 3520 8188
rect 3456 8128 3520 8132
rect 3536 8188 3600 8192
rect 3536 8132 3540 8188
rect 3540 8132 3596 8188
rect 3596 8132 3600 8188
rect 3536 8128 3600 8132
rect 4859 8188 4923 8192
rect 4859 8132 4863 8188
rect 4863 8132 4919 8188
rect 4919 8132 4923 8188
rect 4859 8128 4923 8132
rect 4939 8188 5003 8192
rect 4939 8132 4943 8188
rect 4943 8132 4999 8188
rect 4999 8132 5003 8188
rect 4939 8128 5003 8132
rect 5019 8188 5083 8192
rect 5019 8132 5023 8188
rect 5023 8132 5079 8188
rect 5079 8132 5083 8188
rect 5019 8128 5083 8132
rect 5099 8188 5163 8192
rect 5099 8132 5103 8188
rect 5103 8132 5159 8188
rect 5159 8132 5163 8188
rect 5099 8128 5163 8132
rect 6422 8188 6486 8192
rect 6422 8132 6426 8188
rect 6426 8132 6482 8188
rect 6482 8132 6486 8188
rect 6422 8128 6486 8132
rect 6502 8188 6566 8192
rect 6502 8132 6506 8188
rect 6506 8132 6562 8188
rect 6562 8132 6566 8188
rect 6502 8128 6566 8132
rect 6582 8188 6646 8192
rect 6582 8132 6586 8188
rect 6586 8132 6642 8188
rect 6642 8132 6646 8188
rect 6582 8128 6646 8132
rect 6662 8188 6726 8192
rect 6662 8132 6666 8188
rect 6666 8132 6722 8188
rect 6722 8132 6726 8188
rect 6662 8128 6726 8132
rect 2393 7644 2457 7648
rect 2393 7588 2397 7644
rect 2397 7588 2453 7644
rect 2453 7588 2457 7644
rect 2393 7584 2457 7588
rect 2473 7644 2537 7648
rect 2473 7588 2477 7644
rect 2477 7588 2533 7644
rect 2533 7588 2537 7644
rect 2473 7584 2537 7588
rect 2553 7644 2617 7648
rect 2553 7588 2557 7644
rect 2557 7588 2613 7644
rect 2613 7588 2617 7644
rect 2553 7584 2617 7588
rect 2633 7644 2697 7648
rect 2633 7588 2637 7644
rect 2637 7588 2693 7644
rect 2693 7588 2697 7644
rect 2633 7584 2697 7588
rect 3956 7644 4020 7648
rect 3956 7588 3960 7644
rect 3960 7588 4016 7644
rect 4016 7588 4020 7644
rect 3956 7584 4020 7588
rect 4036 7644 4100 7648
rect 4036 7588 4040 7644
rect 4040 7588 4096 7644
rect 4096 7588 4100 7644
rect 4036 7584 4100 7588
rect 4116 7644 4180 7648
rect 4116 7588 4120 7644
rect 4120 7588 4176 7644
rect 4176 7588 4180 7644
rect 4116 7584 4180 7588
rect 4196 7644 4260 7648
rect 4196 7588 4200 7644
rect 4200 7588 4256 7644
rect 4256 7588 4260 7644
rect 4196 7584 4260 7588
rect 5519 7644 5583 7648
rect 5519 7588 5523 7644
rect 5523 7588 5579 7644
rect 5579 7588 5583 7644
rect 5519 7584 5583 7588
rect 5599 7644 5663 7648
rect 5599 7588 5603 7644
rect 5603 7588 5659 7644
rect 5659 7588 5663 7644
rect 5599 7584 5663 7588
rect 5679 7644 5743 7648
rect 5679 7588 5683 7644
rect 5683 7588 5739 7644
rect 5739 7588 5743 7644
rect 5679 7584 5743 7588
rect 5759 7644 5823 7648
rect 5759 7588 5763 7644
rect 5763 7588 5819 7644
rect 5819 7588 5823 7644
rect 5759 7584 5823 7588
rect 7082 7644 7146 7648
rect 7082 7588 7086 7644
rect 7086 7588 7142 7644
rect 7142 7588 7146 7644
rect 7082 7584 7146 7588
rect 7162 7644 7226 7648
rect 7162 7588 7166 7644
rect 7166 7588 7222 7644
rect 7222 7588 7226 7644
rect 7162 7584 7226 7588
rect 7242 7644 7306 7648
rect 7242 7588 7246 7644
rect 7246 7588 7302 7644
rect 7302 7588 7306 7644
rect 7242 7584 7306 7588
rect 7322 7644 7386 7648
rect 7322 7588 7326 7644
rect 7326 7588 7382 7644
rect 7382 7588 7386 7644
rect 7322 7584 7386 7588
rect 1733 7100 1797 7104
rect 1733 7044 1737 7100
rect 1737 7044 1793 7100
rect 1793 7044 1797 7100
rect 1733 7040 1797 7044
rect 1813 7100 1877 7104
rect 1813 7044 1817 7100
rect 1817 7044 1873 7100
rect 1873 7044 1877 7100
rect 1813 7040 1877 7044
rect 1893 7100 1957 7104
rect 1893 7044 1897 7100
rect 1897 7044 1953 7100
rect 1953 7044 1957 7100
rect 1893 7040 1957 7044
rect 1973 7100 2037 7104
rect 1973 7044 1977 7100
rect 1977 7044 2033 7100
rect 2033 7044 2037 7100
rect 1973 7040 2037 7044
rect 3296 7100 3360 7104
rect 3296 7044 3300 7100
rect 3300 7044 3356 7100
rect 3356 7044 3360 7100
rect 3296 7040 3360 7044
rect 3376 7100 3440 7104
rect 3376 7044 3380 7100
rect 3380 7044 3436 7100
rect 3436 7044 3440 7100
rect 3376 7040 3440 7044
rect 3456 7100 3520 7104
rect 3456 7044 3460 7100
rect 3460 7044 3516 7100
rect 3516 7044 3520 7100
rect 3456 7040 3520 7044
rect 3536 7100 3600 7104
rect 3536 7044 3540 7100
rect 3540 7044 3596 7100
rect 3596 7044 3600 7100
rect 3536 7040 3600 7044
rect 4859 7100 4923 7104
rect 4859 7044 4863 7100
rect 4863 7044 4919 7100
rect 4919 7044 4923 7100
rect 4859 7040 4923 7044
rect 4939 7100 5003 7104
rect 4939 7044 4943 7100
rect 4943 7044 4999 7100
rect 4999 7044 5003 7100
rect 4939 7040 5003 7044
rect 5019 7100 5083 7104
rect 5019 7044 5023 7100
rect 5023 7044 5079 7100
rect 5079 7044 5083 7100
rect 5019 7040 5083 7044
rect 5099 7100 5163 7104
rect 5099 7044 5103 7100
rect 5103 7044 5159 7100
rect 5159 7044 5163 7100
rect 5099 7040 5163 7044
rect 6422 7100 6486 7104
rect 6422 7044 6426 7100
rect 6426 7044 6482 7100
rect 6482 7044 6486 7100
rect 6422 7040 6486 7044
rect 6502 7100 6566 7104
rect 6502 7044 6506 7100
rect 6506 7044 6562 7100
rect 6562 7044 6566 7100
rect 6502 7040 6566 7044
rect 6582 7100 6646 7104
rect 6582 7044 6586 7100
rect 6586 7044 6642 7100
rect 6642 7044 6646 7100
rect 6582 7040 6646 7044
rect 6662 7100 6726 7104
rect 6662 7044 6666 7100
rect 6666 7044 6722 7100
rect 6722 7044 6726 7100
rect 6662 7040 6726 7044
rect 2393 6556 2457 6560
rect 2393 6500 2397 6556
rect 2397 6500 2453 6556
rect 2453 6500 2457 6556
rect 2393 6496 2457 6500
rect 2473 6556 2537 6560
rect 2473 6500 2477 6556
rect 2477 6500 2533 6556
rect 2533 6500 2537 6556
rect 2473 6496 2537 6500
rect 2553 6556 2617 6560
rect 2553 6500 2557 6556
rect 2557 6500 2613 6556
rect 2613 6500 2617 6556
rect 2553 6496 2617 6500
rect 2633 6556 2697 6560
rect 2633 6500 2637 6556
rect 2637 6500 2693 6556
rect 2693 6500 2697 6556
rect 2633 6496 2697 6500
rect 3956 6556 4020 6560
rect 3956 6500 3960 6556
rect 3960 6500 4016 6556
rect 4016 6500 4020 6556
rect 3956 6496 4020 6500
rect 4036 6556 4100 6560
rect 4036 6500 4040 6556
rect 4040 6500 4096 6556
rect 4096 6500 4100 6556
rect 4036 6496 4100 6500
rect 4116 6556 4180 6560
rect 4116 6500 4120 6556
rect 4120 6500 4176 6556
rect 4176 6500 4180 6556
rect 4116 6496 4180 6500
rect 4196 6556 4260 6560
rect 4196 6500 4200 6556
rect 4200 6500 4256 6556
rect 4256 6500 4260 6556
rect 4196 6496 4260 6500
rect 5519 6556 5583 6560
rect 5519 6500 5523 6556
rect 5523 6500 5579 6556
rect 5579 6500 5583 6556
rect 5519 6496 5583 6500
rect 5599 6556 5663 6560
rect 5599 6500 5603 6556
rect 5603 6500 5659 6556
rect 5659 6500 5663 6556
rect 5599 6496 5663 6500
rect 5679 6556 5743 6560
rect 5679 6500 5683 6556
rect 5683 6500 5739 6556
rect 5739 6500 5743 6556
rect 5679 6496 5743 6500
rect 5759 6556 5823 6560
rect 5759 6500 5763 6556
rect 5763 6500 5819 6556
rect 5819 6500 5823 6556
rect 5759 6496 5823 6500
rect 7082 6556 7146 6560
rect 7082 6500 7086 6556
rect 7086 6500 7142 6556
rect 7142 6500 7146 6556
rect 7082 6496 7146 6500
rect 7162 6556 7226 6560
rect 7162 6500 7166 6556
rect 7166 6500 7222 6556
rect 7222 6500 7226 6556
rect 7162 6496 7226 6500
rect 7242 6556 7306 6560
rect 7242 6500 7246 6556
rect 7246 6500 7302 6556
rect 7302 6500 7306 6556
rect 7242 6496 7306 6500
rect 7322 6556 7386 6560
rect 7322 6500 7326 6556
rect 7326 6500 7382 6556
rect 7382 6500 7386 6556
rect 7322 6496 7386 6500
rect 1733 6012 1797 6016
rect 1733 5956 1737 6012
rect 1737 5956 1793 6012
rect 1793 5956 1797 6012
rect 1733 5952 1797 5956
rect 1813 6012 1877 6016
rect 1813 5956 1817 6012
rect 1817 5956 1873 6012
rect 1873 5956 1877 6012
rect 1813 5952 1877 5956
rect 1893 6012 1957 6016
rect 1893 5956 1897 6012
rect 1897 5956 1953 6012
rect 1953 5956 1957 6012
rect 1893 5952 1957 5956
rect 1973 6012 2037 6016
rect 1973 5956 1977 6012
rect 1977 5956 2033 6012
rect 2033 5956 2037 6012
rect 1973 5952 2037 5956
rect 3296 6012 3360 6016
rect 3296 5956 3300 6012
rect 3300 5956 3356 6012
rect 3356 5956 3360 6012
rect 3296 5952 3360 5956
rect 3376 6012 3440 6016
rect 3376 5956 3380 6012
rect 3380 5956 3436 6012
rect 3436 5956 3440 6012
rect 3376 5952 3440 5956
rect 3456 6012 3520 6016
rect 3456 5956 3460 6012
rect 3460 5956 3516 6012
rect 3516 5956 3520 6012
rect 3456 5952 3520 5956
rect 3536 6012 3600 6016
rect 3536 5956 3540 6012
rect 3540 5956 3596 6012
rect 3596 5956 3600 6012
rect 3536 5952 3600 5956
rect 4859 6012 4923 6016
rect 4859 5956 4863 6012
rect 4863 5956 4919 6012
rect 4919 5956 4923 6012
rect 4859 5952 4923 5956
rect 4939 6012 5003 6016
rect 4939 5956 4943 6012
rect 4943 5956 4999 6012
rect 4999 5956 5003 6012
rect 4939 5952 5003 5956
rect 5019 6012 5083 6016
rect 5019 5956 5023 6012
rect 5023 5956 5079 6012
rect 5079 5956 5083 6012
rect 5019 5952 5083 5956
rect 5099 6012 5163 6016
rect 5099 5956 5103 6012
rect 5103 5956 5159 6012
rect 5159 5956 5163 6012
rect 5099 5952 5163 5956
rect 6422 6012 6486 6016
rect 6422 5956 6426 6012
rect 6426 5956 6482 6012
rect 6482 5956 6486 6012
rect 6422 5952 6486 5956
rect 6502 6012 6566 6016
rect 6502 5956 6506 6012
rect 6506 5956 6562 6012
rect 6562 5956 6566 6012
rect 6502 5952 6566 5956
rect 6582 6012 6646 6016
rect 6582 5956 6586 6012
rect 6586 5956 6642 6012
rect 6642 5956 6646 6012
rect 6582 5952 6646 5956
rect 6662 6012 6726 6016
rect 6662 5956 6666 6012
rect 6666 5956 6722 6012
rect 6722 5956 6726 6012
rect 6662 5952 6726 5956
rect 2393 5468 2457 5472
rect 2393 5412 2397 5468
rect 2397 5412 2453 5468
rect 2453 5412 2457 5468
rect 2393 5408 2457 5412
rect 2473 5468 2537 5472
rect 2473 5412 2477 5468
rect 2477 5412 2533 5468
rect 2533 5412 2537 5468
rect 2473 5408 2537 5412
rect 2553 5468 2617 5472
rect 2553 5412 2557 5468
rect 2557 5412 2613 5468
rect 2613 5412 2617 5468
rect 2553 5408 2617 5412
rect 2633 5468 2697 5472
rect 2633 5412 2637 5468
rect 2637 5412 2693 5468
rect 2693 5412 2697 5468
rect 2633 5408 2697 5412
rect 3956 5468 4020 5472
rect 3956 5412 3960 5468
rect 3960 5412 4016 5468
rect 4016 5412 4020 5468
rect 3956 5408 4020 5412
rect 4036 5468 4100 5472
rect 4036 5412 4040 5468
rect 4040 5412 4096 5468
rect 4096 5412 4100 5468
rect 4036 5408 4100 5412
rect 4116 5468 4180 5472
rect 4116 5412 4120 5468
rect 4120 5412 4176 5468
rect 4176 5412 4180 5468
rect 4116 5408 4180 5412
rect 4196 5468 4260 5472
rect 4196 5412 4200 5468
rect 4200 5412 4256 5468
rect 4256 5412 4260 5468
rect 4196 5408 4260 5412
rect 5519 5468 5583 5472
rect 5519 5412 5523 5468
rect 5523 5412 5579 5468
rect 5579 5412 5583 5468
rect 5519 5408 5583 5412
rect 5599 5468 5663 5472
rect 5599 5412 5603 5468
rect 5603 5412 5659 5468
rect 5659 5412 5663 5468
rect 5599 5408 5663 5412
rect 5679 5468 5743 5472
rect 5679 5412 5683 5468
rect 5683 5412 5739 5468
rect 5739 5412 5743 5468
rect 5679 5408 5743 5412
rect 5759 5468 5823 5472
rect 5759 5412 5763 5468
rect 5763 5412 5819 5468
rect 5819 5412 5823 5468
rect 5759 5408 5823 5412
rect 7082 5468 7146 5472
rect 7082 5412 7086 5468
rect 7086 5412 7142 5468
rect 7142 5412 7146 5468
rect 7082 5408 7146 5412
rect 7162 5468 7226 5472
rect 7162 5412 7166 5468
rect 7166 5412 7222 5468
rect 7222 5412 7226 5468
rect 7162 5408 7226 5412
rect 7242 5468 7306 5472
rect 7242 5412 7246 5468
rect 7246 5412 7302 5468
rect 7302 5412 7306 5468
rect 7242 5408 7306 5412
rect 7322 5468 7386 5472
rect 7322 5412 7326 5468
rect 7326 5412 7382 5468
rect 7382 5412 7386 5468
rect 7322 5408 7386 5412
rect 1733 4924 1797 4928
rect 1733 4868 1737 4924
rect 1737 4868 1793 4924
rect 1793 4868 1797 4924
rect 1733 4864 1797 4868
rect 1813 4924 1877 4928
rect 1813 4868 1817 4924
rect 1817 4868 1873 4924
rect 1873 4868 1877 4924
rect 1813 4864 1877 4868
rect 1893 4924 1957 4928
rect 1893 4868 1897 4924
rect 1897 4868 1953 4924
rect 1953 4868 1957 4924
rect 1893 4864 1957 4868
rect 1973 4924 2037 4928
rect 1973 4868 1977 4924
rect 1977 4868 2033 4924
rect 2033 4868 2037 4924
rect 1973 4864 2037 4868
rect 3296 4924 3360 4928
rect 3296 4868 3300 4924
rect 3300 4868 3356 4924
rect 3356 4868 3360 4924
rect 3296 4864 3360 4868
rect 3376 4924 3440 4928
rect 3376 4868 3380 4924
rect 3380 4868 3436 4924
rect 3436 4868 3440 4924
rect 3376 4864 3440 4868
rect 3456 4924 3520 4928
rect 3456 4868 3460 4924
rect 3460 4868 3516 4924
rect 3516 4868 3520 4924
rect 3456 4864 3520 4868
rect 3536 4924 3600 4928
rect 3536 4868 3540 4924
rect 3540 4868 3596 4924
rect 3596 4868 3600 4924
rect 3536 4864 3600 4868
rect 4859 4924 4923 4928
rect 4859 4868 4863 4924
rect 4863 4868 4919 4924
rect 4919 4868 4923 4924
rect 4859 4864 4923 4868
rect 4939 4924 5003 4928
rect 4939 4868 4943 4924
rect 4943 4868 4999 4924
rect 4999 4868 5003 4924
rect 4939 4864 5003 4868
rect 5019 4924 5083 4928
rect 5019 4868 5023 4924
rect 5023 4868 5079 4924
rect 5079 4868 5083 4924
rect 5019 4864 5083 4868
rect 5099 4924 5163 4928
rect 5099 4868 5103 4924
rect 5103 4868 5159 4924
rect 5159 4868 5163 4924
rect 5099 4864 5163 4868
rect 6422 4924 6486 4928
rect 6422 4868 6426 4924
rect 6426 4868 6482 4924
rect 6482 4868 6486 4924
rect 6422 4864 6486 4868
rect 6502 4924 6566 4928
rect 6502 4868 6506 4924
rect 6506 4868 6562 4924
rect 6562 4868 6566 4924
rect 6502 4864 6566 4868
rect 6582 4924 6646 4928
rect 6582 4868 6586 4924
rect 6586 4868 6642 4924
rect 6642 4868 6646 4924
rect 6582 4864 6646 4868
rect 6662 4924 6726 4928
rect 6662 4868 6666 4924
rect 6666 4868 6722 4924
rect 6722 4868 6726 4924
rect 6662 4864 6726 4868
rect 2393 4380 2457 4384
rect 2393 4324 2397 4380
rect 2397 4324 2453 4380
rect 2453 4324 2457 4380
rect 2393 4320 2457 4324
rect 2473 4380 2537 4384
rect 2473 4324 2477 4380
rect 2477 4324 2533 4380
rect 2533 4324 2537 4380
rect 2473 4320 2537 4324
rect 2553 4380 2617 4384
rect 2553 4324 2557 4380
rect 2557 4324 2613 4380
rect 2613 4324 2617 4380
rect 2553 4320 2617 4324
rect 2633 4380 2697 4384
rect 2633 4324 2637 4380
rect 2637 4324 2693 4380
rect 2693 4324 2697 4380
rect 2633 4320 2697 4324
rect 3956 4380 4020 4384
rect 3956 4324 3960 4380
rect 3960 4324 4016 4380
rect 4016 4324 4020 4380
rect 3956 4320 4020 4324
rect 4036 4380 4100 4384
rect 4036 4324 4040 4380
rect 4040 4324 4096 4380
rect 4096 4324 4100 4380
rect 4036 4320 4100 4324
rect 4116 4380 4180 4384
rect 4116 4324 4120 4380
rect 4120 4324 4176 4380
rect 4176 4324 4180 4380
rect 4116 4320 4180 4324
rect 4196 4380 4260 4384
rect 4196 4324 4200 4380
rect 4200 4324 4256 4380
rect 4256 4324 4260 4380
rect 4196 4320 4260 4324
rect 5519 4380 5583 4384
rect 5519 4324 5523 4380
rect 5523 4324 5579 4380
rect 5579 4324 5583 4380
rect 5519 4320 5583 4324
rect 5599 4380 5663 4384
rect 5599 4324 5603 4380
rect 5603 4324 5659 4380
rect 5659 4324 5663 4380
rect 5599 4320 5663 4324
rect 5679 4380 5743 4384
rect 5679 4324 5683 4380
rect 5683 4324 5739 4380
rect 5739 4324 5743 4380
rect 5679 4320 5743 4324
rect 5759 4380 5823 4384
rect 5759 4324 5763 4380
rect 5763 4324 5819 4380
rect 5819 4324 5823 4380
rect 5759 4320 5823 4324
rect 7082 4380 7146 4384
rect 7082 4324 7086 4380
rect 7086 4324 7142 4380
rect 7142 4324 7146 4380
rect 7082 4320 7146 4324
rect 7162 4380 7226 4384
rect 7162 4324 7166 4380
rect 7166 4324 7222 4380
rect 7222 4324 7226 4380
rect 7162 4320 7226 4324
rect 7242 4380 7306 4384
rect 7242 4324 7246 4380
rect 7246 4324 7302 4380
rect 7302 4324 7306 4380
rect 7242 4320 7306 4324
rect 7322 4380 7386 4384
rect 7322 4324 7326 4380
rect 7326 4324 7382 4380
rect 7382 4324 7386 4380
rect 7322 4320 7386 4324
rect 1733 3836 1797 3840
rect 1733 3780 1737 3836
rect 1737 3780 1793 3836
rect 1793 3780 1797 3836
rect 1733 3776 1797 3780
rect 1813 3836 1877 3840
rect 1813 3780 1817 3836
rect 1817 3780 1873 3836
rect 1873 3780 1877 3836
rect 1813 3776 1877 3780
rect 1893 3836 1957 3840
rect 1893 3780 1897 3836
rect 1897 3780 1953 3836
rect 1953 3780 1957 3836
rect 1893 3776 1957 3780
rect 1973 3836 2037 3840
rect 1973 3780 1977 3836
rect 1977 3780 2033 3836
rect 2033 3780 2037 3836
rect 1973 3776 2037 3780
rect 3296 3836 3360 3840
rect 3296 3780 3300 3836
rect 3300 3780 3356 3836
rect 3356 3780 3360 3836
rect 3296 3776 3360 3780
rect 3376 3836 3440 3840
rect 3376 3780 3380 3836
rect 3380 3780 3436 3836
rect 3436 3780 3440 3836
rect 3376 3776 3440 3780
rect 3456 3836 3520 3840
rect 3456 3780 3460 3836
rect 3460 3780 3516 3836
rect 3516 3780 3520 3836
rect 3456 3776 3520 3780
rect 3536 3836 3600 3840
rect 3536 3780 3540 3836
rect 3540 3780 3596 3836
rect 3596 3780 3600 3836
rect 3536 3776 3600 3780
rect 4859 3836 4923 3840
rect 4859 3780 4863 3836
rect 4863 3780 4919 3836
rect 4919 3780 4923 3836
rect 4859 3776 4923 3780
rect 4939 3836 5003 3840
rect 4939 3780 4943 3836
rect 4943 3780 4999 3836
rect 4999 3780 5003 3836
rect 4939 3776 5003 3780
rect 5019 3836 5083 3840
rect 5019 3780 5023 3836
rect 5023 3780 5079 3836
rect 5079 3780 5083 3836
rect 5019 3776 5083 3780
rect 5099 3836 5163 3840
rect 5099 3780 5103 3836
rect 5103 3780 5159 3836
rect 5159 3780 5163 3836
rect 5099 3776 5163 3780
rect 6422 3836 6486 3840
rect 6422 3780 6426 3836
rect 6426 3780 6482 3836
rect 6482 3780 6486 3836
rect 6422 3776 6486 3780
rect 6502 3836 6566 3840
rect 6502 3780 6506 3836
rect 6506 3780 6562 3836
rect 6562 3780 6566 3836
rect 6502 3776 6566 3780
rect 6582 3836 6646 3840
rect 6582 3780 6586 3836
rect 6586 3780 6642 3836
rect 6642 3780 6646 3836
rect 6582 3776 6646 3780
rect 6662 3836 6726 3840
rect 6662 3780 6666 3836
rect 6666 3780 6722 3836
rect 6722 3780 6726 3836
rect 6662 3776 6726 3780
rect 2393 3292 2457 3296
rect 2393 3236 2397 3292
rect 2397 3236 2453 3292
rect 2453 3236 2457 3292
rect 2393 3232 2457 3236
rect 2473 3292 2537 3296
rect 2473 3236 2477 3292
rect 2477 3236 2533 3292
rect 2533 3236 2537 3292
rect 2473 3232 2537 3236
rect 2553 3292 2617 3296
rect 2553 3236 2557 3292
rect 2557 3236 2613 3292
rect 2613 3236 2617 3292
rect 2553 3232 2617 3236
rect 2633 3292 2697 3296
rect 2633 3236 2637 3292
rect 2637 3236 2693 3292
rect 2693 3236 2697 3292
rect 2633 3232 2697 3236
rect 3956 3292 4020 3296
rect 3956 3236 3960 3292
rect 3960 3236 4016 3292
rect 4016 3236 4020 3292
rect 3956 3232 4020 3236
rect 4036 3292 4100 3296
rect 4036 3236 4040 3292
rect 4040 3236 4096 3292
rect 4096 3236 4100 3292
rect 4036 3232 4100 3236
rect 4116 3292 4180 3296
rect 4116 3236 4120 3292
rect 4120 3236 4176 3292
rect 4176 3236 4180 3292
rect 4116 3232 4180 3236
rect 4196 3292 4260 3296
rect 4196 3236 4200 3292
rect 4200 3236 4256 3292
rect 4256 3236 4260 3292
rect 4196 3232 4260 3236
rect 5519 3292 5583 3296
rect 5519 3236 5523 3292
rect 5523 3236 5579 3292
rect 5579 3236 5583 3292
rect 5519 3232 5583 3236
rect 5599 3292 5663 3296
rect 5599 3236 5603 3292
rect 5603 3236 5659 3292
rect 5659 3236 5663 3292
rect 5599 3232 5663 3236
rect 5679 3292 5743 3296
rect 5679 3236 5683 3292
rect 5683 3236 5739 3292
rect 5739 3236 5743 3292
rect 5679 3232 5743 3236
rect 5759 3292 5823 3296
rect 5759 3236 5763 3292
rect 5763 3236 5819 3292
rect 5819 3236 5823 3292
rect 5759 3232 5823 3236
rect 7082 3292 7146 3296
rect 7082 3236 7086 3292
rect 7086 3236 7142 3292
rect 7142 3236 7146 3292
rect 7082 3232 7146 3236
rect 7162 3292 7226 3296
rect 7162 3236 7166 3292
rect 7166 3236 7222 3292
rect 7222 3236 7226 3292
rect 7162 3232 7226 3236
rect 7242 3292 7306 3296
rect 7242 3236 7246 3292
rect 7246 3236 7302 3292
rect 7302 3236 7306 3292
rect 7242 3232 7306 3236
rect 7322 3292 7386 3296
rect 7322 3236 7326 3292
rect 7326 3236 7382 3292
rect 7382 3236 7386 3292
rect 7322 3232 7386 3236
rect 1733 2748 1797 2752
rect 1733 2692 1737 2748
rect 1737 2692 1793 2748
rect 1793 2692 1797 2748
rect 1733 2688 1797 2692
rect 1813 2748 1877 2752
rect 1813 2692 1817 2748
rect 1817 2692 1873 2748
rect 1873 2692 1877 2748
rect 1813 2688 1877 2692
rect 1893 2748 1957 2752
rect 1893 2692 1897 2748
rect 1897 2692 1953 2748
rect 1953 2692 1957 2748
rect 1893 2688 1957 2692
rect 1973 2748 2037 2752
rect 1973 2692 1977 2748
rect 1977 2692 2033 2748
rect 2033 2692 2037 2748
rect 1973 2688 2037 2692
rect 3296 2748 3360 2752
rect 3296 2692 3300 2748
rect 3300 2692 3356 2748
rect 3356 2692 3360 2748
rect 3296 2688 3360 2692
rect 3376 2748 3440 2752
rect 3376 2692 3380 2748
rect 3380 2692 3436 2748
rect 3436 2692 3440 2748
rect 3376 2688 3440 2692
rect 3456 2748 3520 2752
rect 3456 2692 3460 2748
rect 3460 2692 3516 2748
rect 3516 2692 3520 2748
rect 3456 2688 3520 2692
rect 3536 2748 3600 2752
rect 3536 2692 3540 2748
rect 3540 2692 3596 2748
rect 3596 2692 3600 2748
rect 3536 2688 3600 2692
rect 4859 2748 4923 2752
rect 4859 2692 4863 2748
rect 4863 2692 4919 2748
rect 4919 2692 4923 2748
rect 4859 2688 4923 2692
rect 4939 2748 5003 2752
rect 4939 2692 4943 2748
rect 4943 2692 4999 2748
rect 4999 2692 5003 2748
rect 4939 2688 5003 2692
rect 5019 2748 5083 2752
rect 5019 2692 5023 2748
rect 5023 2692 5079 2748
rect 5079 2692 5083 2748
rect 5019 2688 5083 2692
rect 5099 2748 5163 2752
rect 5099 2692 5103 2748
rect 5103 2692 5159 2748
rect 5159 2692 5163 2748
rect 5099 2688 5163 2692
rect 6422 2748 6486 2752
rect 6422 2692 6426 2748
rect 6426 2692 6482 2748
rect 6482 2692 6486 2748
rect 6422 2688 6486 2692
rect 6502 2748 6566 2752
rect 6502 2692 6506 2748
rect 6506 2692 6562 2748
rect 6562 2692 6566 2748
rect 6502 2688 6566 2692
rect 6582 2748 6646 2752
rect 6582 2692 6586 2748
rect 6586 2692 6642 2748
rect 6642 2692 6646 2748
rect 6582 2688 6646 2692
rect 6662 2748 6726 2752
rect 6662 2692 6666 2748
rect 6666 2692 6722 2748
rect 6722 2692 6726 2748
rect 6662 2688 6726 2692
rect 2393 2204 2457 2208
rect 2393 2148 2397 2204
rect 2397 2148 2453 2204
rect 2453 2148 2457 2204
rect 2393 2144 2457 2148
rect 2473 2204 2537 2208
rect 2473 2148 2477 2204
rect 2477 2148 2533 2204
rect 2533 2148 2537 2204
rect 2473 2144 2537 2148
rect 2553 2204 2617 2208
rect 2553 2148 2557 2204
rect 2557 2148 2613 2204
rect 2613 2148 2617 2204
rect 2553 2144 2617 2148
rect 2633 2204 2697 2208
rect 2633 2148 2637 2204
rect 2637 2148 2693 2204
rect 2693 2148 2697 2204
rect 2633 2144 2697 2148
rect 3956 2204 4020 2208
rect 3956 2148 3960 2204
rect 3960 2148 4016 2204
rect 4016 2148 4020 2204
rect 3956 2144 4020 2148
rect 4036 2204 4100 2208
rect 4036 2148 4040 2204
rect 4040 2148 4096 2204
rect 4096 2148 4100 2204
rect 4036 2144 4100 2148
rect 4116 2204 4180 2208
rect 4116 2148 4120 2204
rect 4120 2148 4176 2204
rect 4176 2148 4180 2204
rect 4116 2144 4180 2148
rect 4196 2204 4260 2208
rect 4196 2148 4200 2204
rect 4200 2148 4256 2204
rect 4256 2148 4260 2204
rect 4196 2144 4260 2148
rect 5519 2204 5583 2208
rect 5519 2148 5523 2204
rect 5523 2148 5579 2204
rect 5579 2148 5583 2204
rect 5519 2144 5583 2148
rect 5599 2204 5663 2208
rect 5599 2148 5603 2204
rect 5603 2148 5659 2204
rect 5659 2148 5663 2204
rect 5599 2144 5663 2148
rect 5679 2204 5743 2208
rect 5679 2148 5683 2204
rect 5683 2148 5739 2204
rect 5739 2148 5743 2204
rect 5679 2144 5743 2148
rect 5759 2204 5823 2208
rect 5759 2148 5763 2204
rect 5763 2148 5819 2204
rect 5819 2148 5823 2204
rect 5759 2144 5823 2148
rect 7082 2204 7146 2208
rect 7082 2148 7086 2204
rect 7086 2148 7142 2204
rect 7142 2148 7146 2204
rect 7082 2144 7146 2148
rect 7162 2204 7226 2208
rect 7162 2148 7166 2204
rect 7166 2148 7222 2204
rect 7222 2148 7226 2204
rect 7162 2144 7226 2148
rect 7242 2204 7306 2208
rect 7242 2148 7246 2204
rect 7246 2148 7302 2204
rect 7302 2148 7306 2204
rect 7242 2144 7306 2148
rect 7322 2204 7386 2208
rect 7322 2148 7326 2204
rect 7326 2148 7382 2204
rect 7382 2148 7386 2204
rect 7322 2144 7386 2148
<< metal4 >>
rect 1725 8192 2045 8208
rect 1725 8128 1733 8192
rect 1797 8128 1813 8192
rect 1877 8128 1893 8192
rect 1957 8128 1973 8192
rect 2037 8128 2045 8192
rect 1725 7526 2045 8128
rect 1725 7290 1767 7526
rect 2003 7290 2045 7526
rect 1725 7104 2045 7290
rect 1725 7040 1733 7104
rect 1797 7040 1813 7104
rect 1877 7040 1893 7104
rect 1957 7040 1973 7104
rect 2037 7040 2045 7104
rect 1725 6031 2045 7040
rect 1725 6016 1767 6031
rect 2003 6016 2045 6031
rect 1725 5952 1733 6016
rect 2037 5952 2045 6016
rect 1725 5795 1767 5952
rect 2003 5795 2045 5952
rect 1725 4928 2045 5795
rect 1725 4864 1733 4928
rect 1797 4864 1813 4928
rect 1877 4864 1893 4928
rect 1957 4864 1973 4928
rect 2037 4864 2045 4928
rect 1725 4536 2045 4864
rect 1725 4300 1767 4536
rect 2003 4300 2045 4536
rect 1725 3840 2045 4300
rect 1725 3776 1733 3840
rect 1797 3776 1813 3840
rect 1877 3776 1893 3840
rect 1957 3776 1973 3840
rect 2037 3776 2045 3840
rect 1725 3041 2045 3776
rect 1725 2805 1767 3041
rect 2003 2805 2045 3041
rect 1725 2752 2045 2805
rect 1725 2688 1733 2752
rect 1797 2688 1813 2752
rect 1877 2688 1893 2752
rect 1957 2688 1973 2752
rect 2037 2688 2045 2752
rect 1725 2128 2045 2688
rect 2385 8186 2705 8228
rect 2385 7950 2427 8186
rect 2663 7950 2705 8186
rect 2385 7648 2705 7950
rect 2385 7584 2393 7648
rect 2457 7584 2473 7648
rect 2537 7584 2553 7648
rect 2617 7584 2633 7648
rect 2697 7584 2705 7648
rect 2385 6691 2705 7584
rect 2385 6560 2427 6691
rect 2663 6560 2705 6691
rect 2385 6496 2393 6560
rect 2697 6496 2705 6560
rect 2385 6455 2427 6496
rect 2663 6455 2705 6496
rect 2385 5472 2705 6455
rect 2385 5408 2393 5472
rect 2457 5408 2473 5472
rect 2537 5408 2553 5472
rect 2617 5408 2633 5472
rect 2697 5408 2705 5472
rect 2385 5196 2705 5408
rect 2385 4960 2427 5196
rect 2663 4960 2705 5196
rect 2385 4384 2705 4960
rect 2385 4320 2393 4384
rect 2457 4320 2473 4384
rect 2537 4320 2553 4384
rect 2617 4320 2633 4384
rect 2697 4320 2705 4384
rect 2385 3701 2705 4320
rect 2385 3465 2427 3701
rect 2663 3465 2705 3701
rect 2385 3296 2705 3465
rect 2385 3232 2393 3296
rect 2457 3232 2473 3296
rect 2537 3232 2553 3296
rect 2617 3232 2633 3296
rect 2697 3232 2705 3296
rect 2385 2208 2705 3232
rect 2385 2144 2393 2208
rect 2457 2144 2473 2208
rect 2537 2144 2553 2208
rect 2617 2144 2633 2208
rect 2697 2144 2705 2208
rect 2385 2128 2705 2144
rect 3288 8192 3608 8208
rect 3288 8128 3296 8192
rect 3360 8128 3376 8192
rect 3440 8128 3456 8192
rect 3520 8128 3536 8192
rect 3600 8128 3608 8192
rect 3288 7526 3608 8128
rect 3288 7290 3330 7526
rect 3566 7290 3608 7526
rect 3288 7104 3608 7290
rect 3288 7040 3296 7104
rect 3360 7040 3376 7104
rect 3440 7040 3456 7104
rect 3520 7040 3536 7104
rect 3600 7040 3608 7104
rect 3288 6031 3608 7040
rect 3288 6016 3330 6031
rect 3566 6016 3608 6031
rect 3288 5952 3296 6016
rect 3600 5952 3608 6016
rect 3288 5795 3330 5952
rect 3566 5795 3608 5952
rect 3288 4928 3608 5795
rect 3288 4864 3296 4928
rect 3360 4864 3376 4928
rect 3440 4864 3456 4928
rect 3520 4864 3536 4928
rect 3600 4864 3608 4928
rect 3288 4536 3608 4864
rect 3288 4300 3330 4536
rect 3566 4300 3608 4536
rect 3288 3840 3608 4300
rect 3288 3776 3296 3840
rect 3360 3776 3376 3840
rect 3440 3776 3456 3840
rect 3520 3776 3536 3840
rect 3600 3776 3608 3840
rect 3288 3041 3608 3776
rect 3288 2805 3330 3041
rect 3566 2805 3608 3041
rect 3288 2752 3608 2805
rect 3288 2688 3296 2752
rect 3360 2688 3376 2752
rect 3440 2688 3456 2752
rect 3520 2688 3536 2752
rect 3600 2688 3608 2752
rect 3288 2128 3608 2688
rect 3948 8186 4268 8228
rect 3948 7950 3990 8186
rect 4226 7950 4268 8186
rect 3948 7648 4268 7950
rect 3948 7584 3956 7648
rect 4020 7584 4036 7648
rect 4100 7584 4116 7648
rect 4180 7584 4196 7648
rect 4260 7584 4268 7648
rect 3948 6691 4268 7584
rect 3948 6560 3990 6691
rect 4226 6560 4268 6691
rect 3948 6496 3956 6560
rect 4260 6496 4268 6560
rect 3948 6455 3990 6496
rect 4226 6455 4268 6496
rect 3948 5472 4268 6455
rect 3948 5408 3956 5472
rect 4020 5408 4036 5472
rect 4100 5408 4116 5472
rect 4180 5408 4196 5472
rect 4260 5408 4268 5472
rect 3948 5196 4268 5408
rect 3948 4960 3990 5196
rect 4226 4960 4268 5196
rect 3948 4384 4268 4960
rect 3948 4320 3956 4384
rect 4020 4320 4036 4384
rect 4100 4320 4116 4384
rect 4180 4320 4196 4384
rect 4260 4320 4268 4384
rect 3948 3701 4268 4320
rect 3948 3465 3990 3701
rect 4226 3465 4268 3701
rect 3948 3296 4268 3465
rect 3948 3232 3956 3296
rect 4020 3232 4036 3296
rect 4100 3232 4116 3296
rect 4180 3232 4196 3296
rect 4260 3232 4268 3296
rect 3948 2208 4268 3232
rect 3948 2144 3956 2208
rect 4020 2144 4036 2208
rect 4100 2144 4116 2208
rect 4180 2144 4196 2208
rect 4260 2144 4268 2208
rect 3948 2128 4268 2144
rect 4851 8192 5171 8208
rect 4851 8128 4859 8192
rect 4923 8128 4939 8192
rect 5003 8128 5019 8192
rect 5083 8128 5099 8192
rect 5163 8128 5171 8192
rect 4851 7526 5171 8128
rect 4851 7290 4893 7526
rect 5129 7290 5171 7526
rect 4851 7104 5171 7290
rect 4851 7040 4859 7104
rect 4923 7040 4939 7104
rect 5003 7040 5019 7104
rect 5083 7040 5099 7104
rect 5163 7040 5171 7104
rect 4851 6031 5171 7040
rect 4851 6016 4893 6031
rect 5129 6016 5171 6031
rect 4851 5952 4859 6016
rect 5163 5952 5171 6016
rect 4851 5795 4893 5952
rect 5129 5795 5171 5952
rect 4851 4928 5171 5795
rect 4851 4864 4859 4928
rect 4923 4864 4939 4928
rect 5003 4864 5019 4928
rect 5083 4864 5099 4928
rect 5163 4864 5171 4928
rect 4851 4536 5171 4864
rect 4851 4300 4893 4536
rect 5129 4300 5171 4536
rect 4851 3840 5171 4300
rect 4851 3776 4859 3840
rect 4923 3776 4939 3840
rect 5003 3776 5019 3840
rect 5083 3776 5099 3840
rect 5163 3776 5171 3840
rect 4851 3041 5171 3776
rect 4851 2805 4893 3041
rect 5129 2805 5171 3041
rect 4851 2752 5171 2805
rect 4851 2688 4859 2752
rect 4923 2688 4939 2752
rect 5003 2688 5019 2752
rect 5083 2688 5099 2752
rect 5163 2688 5171 2752
rect 4851 2128 5171 2688
rect 5511 8186 5831 8228
rect 5511 7950 5553 8186
rect 5789 7950 5831 8186
rect 5511 7648 5831 7950
rect 5511 7584 5519 7648
rect 5583 7584 5599 7648
rect 5663 7584 5679 7648
rect 5743 7584 5759 7648
rect 5823 7584 5831 7648
rect 5511 6691 5831 7584
rect 5511 6560 5553 6691
rect 5789 6560 5831 6691
rect 5511 6496 5519 6560
rect 5823 6496 5831 6560
rect 5511 6455 5553 6496
rect 5789 6455 5831 6496
rect 5511 5472 5831 6455
rect 5511 5408 5519 5472
rect 5583 5408 5599 5472
rect 5663 5408 5679 5472
rect 5743 5408 5759 5472
rect 5823 5408 5831 5472
rect 5511 5196 5831 5408
rect 5511 4960 5553 5196
rect 5789 4960 5831 5196
rect 5511 4384 5831 4960
rect 5511 4320 5519 4384
rect 5583 4320 5599 4384
rect 5663 4320 5679 4384
rect 5743 4320 5759 4384
rect 5823 4320 5831 4384
rect 5511 3701 5831 4320
rect 5511 3465 5553 3701
rect 5789 3465 5831 3701
rect 5511 3296 5831 3465
rect 5511 3232 5519 3296
rect 5583 3232 5599 3296
rect 5663 3232 5679 3296
rect 5743 3232 5759 3296
rect 5823 3232 5831 3296
rect 5511 2208 5831 3232
rect 5511 2144 5519 2208
rect 5583 2144 5599 2208
rect 5663 2144 5679 2208
rect 5743 2144 5759 2208
rect 5823 2144 5831 2208
rect 5511 2128 5831 2144
rect 6414 8192 6734 8208
rect 6414 8128 6422 8192
rect 6486 8128 6502 8192
rect 6566 8128 6582 8192
rect 6646 8128 6662 8192
rect 6726 8128 6734 8192
rect 6414 7526 6734 8128
rect 6414 7290 6456 7526
rect 6692 7290 6734 7526
rect 6414 7104 6734 7290
rect 6414 7040 6422 7104
rect 6486 7040 6502 7104
rect 6566 7040 6582 7104
rect 6646 7040 6662 7104
rect 6726 7040 6734 7104
rect 6414 6031 6734 7040
rect 6414 6016 6456 6031
rect 6692 6016 6734 6031
rect 6414 5952 6422 6016
rect 6726 5952 6734 6016
rect 6414 5795 6456 5952
rect 6692 5795 6734 5952
rect 6414 4928 6734 5795
rect 6414 4864 6422 4928
rect 6486 4864 6502 4928
rect 6566 4864 6582 4928
rect 6646 4864 6662 4928
rect 6726 4864 6734 4928
rect 6414 4536 6734 4864
rect 6414 4300 6456 4536
rect 6692 4300 6734 4536
rect 6414 3840 6734 4300
rect 6414 3776 6422 3840
rect 6486 3776 6502 3840
rect 6566 3776 6582 3840
rect 6646 3776 6662 3840
rect 6726 3776 6734 3840
rect 6414 3041 6734 3776
rect 6414 2805 6456 3041
rect 6692 2805 6734 3041
rect 6414 2752 6734 2805
rect 6414 2688 6422 2752
rect 6486 2688 6502 2752
rect 6566 2688 6582 2752
rect 6646 2688 6662 2752
rect 6726 2688 6734 2752
rect 6414 2128 6734 2688
rect 7074 8186 7394 8228
rect 7074 7950 7116 8186
rect 7352 7950 7394 8186
rect 7074 7648 7394 7950
rect 7074 7584 7082 7648
rect 7146 7584 7162 7648
rect 7226 7584 7242 7648
rect 7306 7584 7322 7648
rect 7386 7584 7394 7648
rect 7074 6691 7394 7584
rect 7074 6560 7116 6691
rect 7352 6560 7394 6691
rect 7074 6496 7082 6560
rect 7386 6496 7394 6560
rect 7074 6455 7116 6496
rect 7352 6455 7394 6496
rect 7074 5472 7394 6455
rect 7074 5408 7082 5472
rect 7146 5408 7162 5472
rect 7226 5408 7242 5472
rect 7306 5408 7322 5472
rect 7386 5408 7394 5472
rect 7074 5196 7394 5408
rect 7074 4960 7116 5196
rect 7352 4960 7394 5196
rect 7074 4384 7394 4960
rect 7074 4320 7082 4384
rect 7146 4320 7162 4384
rect 7226 4320 7242 4384
rect 7306 4320 7322 4384
rect 7386 4320 7394 4384
rect 7074 3701 7394 4320
rect 7074 3465 7116 3701
rect 7352 3465 7394 3701
rect 7074 3296 7394 3465
rect 7074 3232 7082 3296
rect 7146 3232 7162 3296
rect 7226 3232 7242 3296
rect 7306 3232 7322 3296
rect 7386 3232 7394 3296
rect 7074 2208 7394 3232
rect 7074 2144 7082 2208
rect 7146 2144 7162 2208
rect 7226 2144 7242 2208
rect 7306 2144 7322 2208
rect 7386 2144 7394 2208
rect 7074 2128 7394 2144
<< via4 >>
rect 1767 7290 2003 7526
rect 1767 6016 2003 6031
rect 1767 5952 1797 6016
rect 1797 5952 1813 6016
rect 1813 5952 1877 6016
rect 1877 5952 1893 6016
rect 1893 5952 1957 6016
rect 1957 5952 1973 6016
rect 1973 5952 2003 6016
rect 1767 5795 2003 5952
rect 1767 4300 2003 4536
rect 1767 2805 2003 3041
rect 2427 7950 2663 8186
rect 2427 6560 2663 6691
rect 2427 6496 2457 6560
rect 2457 6496 2473 6560
rect 2473 6496 2537 6560
rect 2537 6496 2553 6560
rect 2553 6496 2617 6560
rect 2617 6496 2633 6560
rect 2633 6496 2663 6560
rect 2427 6455 2663 6496
rect 2427 4960 2663 5196
rect 2427 3465 2663 3701
rect 3330 7290 3566 7526
rect 3330 6016 3566 6031
rect 3330 5952 3360 6016
rect 3360 5952 3376 6016
rect 3376 5952 3440 6016
rect 3440 5952 3456 6016
rect 3456 5952 3520 6016
rect 3520 5952 3536 6016
rect 3536 5952 3566 6016
rect 3330 5795 3566 5952
rect 3330 4300 3566 4536
rect 3330 2805 3566 3041
rect 3990 7950 4226 8186
rect 3990 6560 4226 6691
rect 3990 6496 4020 6560
rect 4020 6496 4036 6560
rect 4036 6496 4100 6560
rect 4100 6496 4116 6560
rect 4116 6496 4180 6560
rect 4180 6496 4196 6560
rect 4196 6496 4226 6560
rect 3990 6455 4226 6496
rect 3990 4960 4226 5196
rect 3990 3465 4226 3701
rect 4893 7290 5129 7526
rect 4893 6016 5129 6031
rect 4893 5952 4923 6016
rect 4923 5952 4939 6016
rect 4939 5952 5003 6016
rect 5003 5952 5019 6016
rect 5019 5952 5083 6016
rect 5083 5952 5099 6016
rect 5099 5952 5129 6016
rect 4893 5795 5129 5952
rect 4893 4300 5129 4536
rect 4893 2805 5129 3041
rect 5553 7950 5789 8186
rect 5553 6560 5789 6691
rect 5553 6496 5583 6560
rect 5583 6496 5599 6560
rect 5599 6496 5663 6560
rect 5663 6496 5679 6560
rect 5679 6496 5743 6560
rect 5743 6496 5759 6560
rect 5759 6496 5789 6560
rect 5553 6455 5789 6496
rect 5553 4960 5789 5196
rect 5553 3465 5789 3701
rect 6456 7290 6692 7526
rect 6456 6016 6692 6031
rect 6456 5952 6486 6016
rect 6486 5952 6502 6016
rect 6502 5952 6566 6016
rect 6566 5952 6582 6016
rect 6582 5952 6646 6016
rect 6646 5952 6662 6016
rect 6662 5952 6692 6016
rect 6456 5795 6692 5952
rect 6456 4300 6692 4536
rect 6456 2805 6692 3041
rect 7116 7950 7352 8186
rect 7116 6560 7352 6691
rect 7116 6496 7146 6560
rect 7146 6496 7162 6560
rect 7162 6496 7226 6560
rect 7226 6496 7242 6560
rect 7242 6496 7306 6560
rect 7306 6496 7322 6560
rect 7322 6496 7352 6560
rect 7116 6455 7352 6496
rect 7116 4960 7352 5196
rect 7116 3465 7352 3701
<< metal5 >>
rect 1056 8186 7408 8228
rect 1056 7950 2427 8186
rect 2663 7950 3990 8186
rect 4226 7950 5553 8186
rect 5789 7950 7116 8186
rect 7352 7950 7408 8186
rect 1056 7908 7408 7950
rect 1056 7526 7408 7568
rect 1056 7290 1767 7526
rect 2003 7290 3330 7526
rect 3566 7290 4893 7526
rect 5129 7290 6456 7526
rect 6692 7290 7408 7526
rect 1056 7248 7408 7290
rect 1056 6691 7408 6733
rect 1056 6455 2427 6691
rect 2663 6455 3990 6691
rect 4226 6455 5553 6691
rect 5789 6455 7116 6691
rect 7352 6455 7408 6691
rect 1056 6413 7408 6455
rect 1056 6031 7408 6073
rect 1056 5795 1767 6031
rect 2003 5795 3330 6031
rect 3566 5795 4893 6031
rect 5129 5795 6456 6031
rect 6692 5795 7408 6031
rect 1056 5753 7408 5795
rect 1056 5196 7408 5238
rect 1056 4960 2427 5196
rect 2663 4960 3990 5196
rect 4226 4960 5553 5196
rect 5789 4960 7116 5196
rect 7352 4960 7408 5196
rect 1056 4918 7408 4960
rect 1056 4536 7408 4578
rect 1056 4300 1767 4536
rect 2003 4300 3330 4536
rect 3566 4300 4893 4536
rect 5129 4300 6456 4536
rect 6692 4300 7408 4536
rect 1056 4258 7408 4300
rect 1056 3701 7408 3743
rect 1056 3465 2427 3701
rect 2663 3465 3990 3701
rect 4226 3465 5553 3701
rect 5789 3465 7116 3701
rect 7352 3465 7408 3701
rect 1056 3423 7408 3465
rect 1056 3041 7408 3083
rect 1056 2805 1767 3041
rect 2003 2805 3330 3041
rect 3566 2805 4893 3041
rect 5129 2805 6456 3041
rect 6692 2805 7408 3041
rect 1056 2763 7408 2805
use sky130_fd_sc_hd__xnor2_1  _2_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5152 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _3_
timestamp 1704896540
transform 1 0 3864 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _4_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _5_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1704896540
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1704896540
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_35
timestamp 1704896540
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_47
timestamp 1704896540
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_7
timestamp 1704896540
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_19
timestamp 1704896540
transform 1 0 2852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_23
timestamp 1704896540
transform 1 0 3220 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_44
timestamp 1704896540
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 1704896540
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1704896540
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1704896540
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1704896540
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_57
timestamp 1704896540
transform 1 0 6348 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform -1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1704896540
transform 1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_11
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_12
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_13
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_14
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_15
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_16
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_17
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_18
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_19
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_20
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_21
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 7360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_24
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_25
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_26
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_27
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_28
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_30
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_31
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_32
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_33
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_34
timestamp 1704896540
transform 1 0 6256 0 1 7616
box -38 -48 130 592
<< labels >>
flabel metal4 s 2385 2128 2705 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3948 2128 4268 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5511 2128 5831 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7074 2128 7394 8228 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3423 7408 3743 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4918 7408 5238 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6413 7408 6733 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7908 7408 8228 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1725 2128 2045 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3288 2128 3608 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4851 2128 5171 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6414 2128 6734 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2763 7408 3083 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4258 7408 4578 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5753 7408 6073 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7248 7408 7568 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 a
port 2 nsew signal input
flabel metal3 s 7735 4768 8535 4888 0 FreeSans 480 0 0 0 b
port 3 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 cin
port 4 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 co
port 5 nsew signal output
flabel metal3 s 7735 5448 8535 5568 0 FreeSans 480 0 0 0 s
port 6 nsew signal output
rlabel via1 4249 7616 4249 7616 0 VGND
rlabel metal1 4232 8160 4232 8160 0 VPWR
rlabel metal1 4002 5100 4002 5100 0 _0_
rlabel metal2 4002 4794 4002 4794 0 _1_
rlabel metal3 1050 5508 1050 5508 0 a
rlabel metal2 7038 5015 7038 5015 0 b
rlabel metal3 751 4148 751 4148 0 cin
rlabel metal3 751 4828 751 4828 0 co
rlabel metal2 3358 5372 3358 5372 0 net1
rlabel metal1 4922 5134 4922 5134 0 net2
rlabel metal1 3634 5168 3634 5168 0 net3
rlabel metal1 3496 4794 3496 4794 0 net4
rlabel metal1 5612 5338 5612 5338 0 net5
rlabel metal1 7222 5542 7222 5542 0 s
<< properties >>
string FIXED_BBOX 0 0 8535 10679
<< end >>
